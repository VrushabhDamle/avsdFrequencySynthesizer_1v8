*PLL
.include sky130nm.lib
.option scale = 0.01u
xx1 Clk_Ref Clk_Out_by_8 up down pd
xx2 up down VCtrl cp

*Loop Filter
r1 VCtrl rc1 490
c1 rc1 0 215f
r2 rc1 rc2 490
c2 rc2 0 210f
r3 rc2 rc3 490
c3 rc3 0 205f

xx3 rc3 Clk_Out vco

xx4 Clk_Out Clk_Out_by_2 fd
xx5 Clk_Out_by_2 Clk_Out_by_4 fd
xx6 Clk_Out_by_4 Clk_Out_by_8 fd

v1 Clk_Ref 0 PULSE 0 1.8 0 6ps 6ps 0.333us 0.666us

.ic v(VCtrl) = 0
.ic v(Clk_Out_by_2) = 0
.ic v(Clk_Out_by_4) = 1.8
.ic v(Clk_Out_by_8) = 0
.control
tran 0.1ns 200us
*plot v(Clk_Ref) v(Clk_Out_by_8) v(Clk_Out_by_4)+2 v(Clk_Out_by_2)+4 v(Clk_Out)+6 v(up)+8 v(down)+10 v(VCtrl)+12
*plot v(Clk_Ref) v(Clk_Out_by_8)+2 v(Clk_Out)+4
plot v(Clk_Out)
.endc

*PFD
.subckt pd Clk_Ref Clk2 Up Down 
XM1000 VDD a_7_412# a_460_368# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=1664.03 pd=142.146 as=2232 ps=206
XM1001 GND a_7_412# a_460_368# GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=842.4 pd=91.8 as=1116 ps=134
XM1002 a_264_92# Clk2 a_208_92# GND sky130_fd_pr__nfet_01v8 w=240 l=15
+  ad=7920 pd=546 as=5314.29 ps=321.143
XM1003 VDD Clk2 a_208_92# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=1502.25 pd=128.326 as=2145 ps=196
XM1004 Up a_460_368# GND GND sky130_fd_pr__nfet_01v8 w=48 l=15
+  ad=1392 pd=154 as=1123.2 ps=122.4
XM1005 GND a_264_92# a_485_83# GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=842.4 pd=91.8 as=1116 ps=134
XM1006 a_151_92# Clk_Ref GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=74 as=842.4 ps=91.8
XM1007 VDD a_264_92# a_485_83# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=1664.03 pd=142.146 as=2232 ps=206
XM1008 Down a_485_83# VDD VDD sky130_fd_pr__pfet_01v8 w=96 l=15
+  ad=2880 pd=252 as=2218.71 ps=189.528
XM1009 a_7_412# Clk_Ref a_7_356# GND sky130_fd_pr__nfet_01v8 w=240 l=15
+  ad=7920 pd=546 as=5314.29 ps=321.143
XM1010 Up a_460_368# VDD VDD sky130_fd_pr__pfet_01v8 w=96 l=15
+  ad=2880 pd=252 as=2218.71 ps=189.528
XM1011 VDD Clk_Ref a_7_356# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=1502.25 pd=128.326 as=2145 ps=196
XM1012 Down a_485_83# GND GND sky130_fd_pr__nfet_01v8 w=48 l=15
+  ad=1392 pd=154 as=1123.2 ps=122.4
XM1013 Clk_Ref Clk_Ref a_7_412# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=2145 pd=196 as=2145 ps=196
XM1014 a_7_299# Clk2 GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=74 as=842.4 ps=91.8
XM1015 a_208_92# Clk2 a_151_92# GND sky130_fd_pr__nfet_01v8 w=180 l=15
+  ad=3985.71 pd=240.857 as=5220 ps=370
XM1016 Clk2 Clk2 a_264_92# VDD sky130_fd_pr__pfet_01v8 w=65 l=15
+  ad=2145 pd=196 as=2145 ps=196
XM1017 a_7_356# Clk_Ref a_7_299# GND sky130_fd_pr__nfet_01v8 w=180 l=15
+  ad=3985.71 pd=240.857 as=5220 ps=370
C0 Down Up 0.00fF
C1 a_264_92# VDD 0.13fF
C2 a_208_92# a_485_83# 0.02fF
C3 a_460_368# Clk_Ref 0.00fF
C4 Clk2 a_485_83# 0.06fF
C5 a_7_412# VDD 0.14fF
C6 Up VDD 0.13fF
C7 a_460_368# a_485_83# 0.01fF
C8 Down VDD 0.56fF
C9 a_264_92# a_208_92# 0.49fF
C10 a_264_92# Clk2 0.27fF
C11 a_264_92# Clk_Ref 0.01fF
C12 a_7_412# a_208_92# 0.01fF
C13 a_7_412# Clk2 0.01fF
C14 a_7_412# Clk_Ref 0.19fF
C15 a_264_92# a_460_368# 0.00fF
C16 a_7_412# a_7_356# 0.49fF
C17 a_264_92# a_485_83# 0.37fF
C18 a_7_412# a_460_368# 0.34fF
C19 Down Clk2 0.02fF
C20 a_7_412# a_485_83# 0.00fF
C21 a_460_368# Up 0.16fF
C22 Up a_485_83# 0.00fF
C23 a_208_92# VDD 0.27fF
C24 Clk2 VDD 0.08fF
C25 VDD Clk_Ref 0.20fF
C26 Down a_485_83# 0.16fF
C27 a_7_356# VDD 0.15fF
C28 a_7_412# a_264_92# 0.03fF
C29 a_460_368# VDD 0.20fF
C30 VDD a_485_83# 0.31fF
C31 a_208_92# Clk2 0.05fF
C32 a_208_92# Clk_Ref 0.01fF
C33 a_7_412# Up 0.01fF
C34 Clk2 Clk_Ref 0.11fF
C35 Down a_264_92# 0.01fF
C36 a_7_356# a_208_92# 0.02fF
C37 a_7_356# Clk2 0.01fF
C38 a_7_356# Clk_Ref 0.10fF
C39 Up GND 0.22fF
C40 VDD GND 4.13fF
C41 a_485_83# GND 0.34fF
C42 a_264_92# GND 0.52fF
C43 a_208_92# GND 0.10fF
C44 a_7_356# GND 0.34fF
C45 a_460_368# GND 0.34fF
C46 a_7_412# GND 0.65fF


*output cap
*c1 up 0 6f
*c2 down 0 6f

v1 VDD GND 1.8
.ends pd


*CP
.subckt cp Up Down Out
XM1000 a_174_531# a_127_486# a_248_475# VDD sky130_fd_pr__pfet_01v8 w=1800 l=15
+  ad=59400 pd=3728.85 as=47294.2 ps=2895.72
XM1001 GND a_340_202# a_462_191# GND sky130_fd_pr__nfet_01v8 w=480 l=15
+  ad=15785.8 pd=1205.27 as=10416.3 ps=592.994
XM1002 a_248_475# a_134_73# Out VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1103.53 pd=67.5667 as=1386 ps=150
XM1003 a_134_73# Down GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1188 pd=138 as=1183.94 ps=90.395
XM1004 VDD ENb a_31_494# VDD sky130_fd_pr__pfet_01v8 w=60 l=15
+  ad=2023.9 pd=185.854 as=2340 ps=198
XM1005 a_248_475# Down a_248_427# VDD sky130_fd_pr__pfet_01v8 w=540 l=15
+  ad=14188.3 pd=868.715 as=17820 ps=1146
XM1006 a_258_74# Up GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1188 pd=138 as=1183.94 ps=90.395
XM1007 GND a_340_202# a_340_202# GND sky130_fd_pr__nfet_01v8 w=44 l=15
+  ad=1447.03 pd=110.483 as=1452 ps=154
XM1008 a_462_143# a_462_143# VDD VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1386 pd=150 as=1416.73 ps=130.098
XM1009 a_174_531# a_127_486# a_127_486# VDD sky130_fd_pr__pfet_01v8 w=44 l=15
+  ad=1452 pd=91.1497 as=1452 ps=154
XM1010 Out Up a_462_191# GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1386 pd=150 as=911.424 ps=51.887
XM1011 a_248_427# a_248_427# GND GND sky130_fd_pr__nfet_01v8 w=42 l=15
+  ad=1386 pd=150 as=1381.26 ps=105.461
XM1012 a_462_191# a_258_74# a_462_143# GND sky130_fd_pr__nfet_01v8 w=540 l=15
+  ad=11718.3 pd=667.119 as=17820 ps=1146
XM1013 a_258_74# Up VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2376 pd=210 as=2428.68 ps=223.024
XM1014 a_134_73# Down VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2376 pd=210 as=2428.68 ps=223.024
C0 a_258_74# VDD 0.18fF
C1 VDD Up 0.21fF
C2 a_248_427# Out 0.00fF
C3 a_258_74# Up 0.09fF
C4 a_462_191# a_340_202# 0.01fF
C5 a_134_73# Down 0.12fF
C6 Down ENb 0.00fF
C7 a_462_191# a_462_143# 0.72fF
C8 a_134_73# VDD 0.16fF
C9 a_248_475# a_248_427# 0.58fF
C10 VDD ENb 0.01fF
C11 a_174_531# a_248_427# 0.25fF
C12 a_134_73# a_258_74# 0.05fF
C13 a_134_73# Up 0.41fF
C14 VDD Out 1.29fF
C15 a_462_191# a_248_427# 0.02fF
C16 a_127_486# Down 0.03fF
C17 a_462_143# a_248_427# 0.01fF
C18 Out Up 0.03fF
C19 a_127_486# VDD 0.05fF
C20 a_174_531# Down 0.02fF
C21 a_248_475# VDD 1.18fF
C22 a_174_531# VDD 2.61fF
C23 a_340_202# VDD 0.02fF
C24 a_340_202# a_258_74# 0.13fF
C25 a_340_202# Up 0.02fF
C26 a_462_191# VDD 0.13fF
C27 a_134_73# Out 0.05fF
C28 a_174_531# a_31_494# 0.12fF
C29 a_462_143# VDD 0.23fF
C30 a_462_191# a_258_74# 0.00fF
C31 a_462_191# Up 0.09fF
C32 a_258_74# a_462_143# 0.02fF
C33 a_462_143# Up 0.08fF
C34 a_127_486# ENb 0.01fF
C35 a_248_427# Down 0.00fF
C36 a_134_73# a_248_475# 0.02fF
C37 a_248_427# VDD 0.14fF
C38 a_134_73# a_174_531# 0.01fF
C39 a_134_73# a_340_202# 0.00fF
C40 a_174_531# ENb 0.01fF
C41 a_258_74# a_248_427# 0.00fF
C42 a_248_475# Out 0.40fF
C43 a_174_531# Out 0.24fF
C44 a_127_486# a_248_475# 0.02fF
C45 a_462_191# Out 0.04fF
C46 a_127_486# a_174_531# 0.13fF
C47 Down VDD 0.05fF
C48 a_462_143# Out 0.02fF
C49 a_134_73# a_248_427# 0.09fF
C50 a_258_74# Down 0.00fF
C51 Down Up 0.15fF
C52 a_174_531# a_248_475# 2.05fF
C53 Up GND 1.42fF
C54 Out GND 2.98fF
C55 VDD GND 0.08fF
C56 a_462_143# GND 0.58fF
C57 a_462_191# GND 0.58fF
C58 a_340_202# GND 0.31fF
C59 a_258_74# GND 0.51fF
C60 a_134_73# GND 2.42fF
C61 a_248_427# GND 0.69fF
C62 a_248_475# GND 0.49fF
C63 a_127_486# GND 0.24fF
C64 a_174_531# GND 1.49fF

*r1 out rc 200
*c1 rc 0 8f

v2 ENb 0 0
v1 VDD GND 1.8
.ends cp


*VCO
.subckt vco in out

X0 a_n29_n330# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X1 a_115_n174# a_15_n174# a_n29_n330# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X2 a_n29_379# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X3 a_515_n174# a_415_n174# a_n29_n730# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X4 a_n29_n630# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X5 out a_n29_n49# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=420 l=15
X6 out a_n29_n49# gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X7 a_215_n174# a_115_n174# a_n29_379# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X8 a_n29_679# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X9 a_315_n174# a_215_n174# a_n29_479# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X10 a_15_n174# a_n29_n49# a_n29_n230# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X11 a_415_n174# a_315_n174# a_n29_n630# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X12 a_n29_n230# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X13 a_n29_279# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X14 a_n29_n530# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X15 a_n29_579# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X16 a_n29_n830# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X17 a_415_n174# a_315_n174# a_n29_579# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X18 a_315_n174# a_215_n174# a_n29_n530# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X19 a_n29_0# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X20 a_515_n174# a_415_n174# a_n29_679# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X21 a_n29_n430# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X22 a_n29_479# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X23 a_215_n174# a_115_n174# a_n29_n430# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X24 a_n29_n730# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X25 a_n29_n49# a_515_n174# a_n29_n830# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X26 a_n29_779# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X27 a_n29_n49# a_515_n174# a_n29_779# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X28 a_n124_86# in gnd SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X29 a_n124_86# a_n124_86# vdd w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=500 l=15
X30 a_15_n174# a_n29_n49# a_n29_0# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15
X31 a_115_n174# a_15_n174# a_n29_279# w_n171_117# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=108 l=15

C0 a_515_n174# a_n29_n630# 0.03fF
C1 a_n29_0# a_n29_n49# 0.04fF
C2 a_n29_n430# a_n124_86# 0.01fF
C3 a_15_n174# gnd 0.01fF
C4 a_n29_479# a_n29_679# 0.14fF
C5 a_n29_n730# out 0.06fF
C6 gnd out 0.14fF
C7 a_n29_n630# a_n29_n230# 0.09fF
C8 a_515_n174# out 0.07fF
C9 a_n29_579# a_n29_n630# 0.01fF
C10 a_115_n174# vdd 0.03fF
C11 a_n29_279# a_n29_579# 0.07fF
C12 a_415_n174# a_n29_n530# 0.03fF
C13 a_n29_n730# a_n29_n49# 0.03fF
C14 a_n29_n49# gnd 0.00fF
C15 a_n29_n630# a_n29_n830# 0.12fF
C16 a_15_n174# a_n29_n230# 0.16fF
C17 a_n29_379# a_n29_679# 0.03fF
C18 a_515_n174# a_n29_n49# 0.37fF
C19 a_n124_86# a_n29_n530# 0.01fF
C20 a_115_n174# a_315_n174# 0.06fF
C21 a_n29_n330# a_115_n174# 0.14fF
C22 a_n29_n430# a_n29_379# 0.01fF
C23 a_415_n174# a_n124_86# 0.00fF
C24 a_n29_n330# in 0.03fF
C25 a_n29_n830# out 0.10fF
C26 a_n29_n230# a_n29_n49# 0.03fF
C27 a_415_n174# w_n171_117# 0.00fF
C28 a_n29_479# a_n29_n530# 0.01fF
C29 a_n29_579# a_n29_n49# 0.01fF
C30 a_n29_279# vdd 1.56fF
C31 a_n124_86# w_n171_117# 0.00fF
C32 a_n29_n830# a_n29_n49# 0.13fF
C33 a_415_n174# a_n29_479# 0.03fF
C34 a_15_n174# vdd 0.03fF
C35 a_n29_n630# a_315_n174# 0.13fF
C36 a_n29_679# a_n29_779# 0.82fF
C37 a_n29_279# a_315_n174# 0.00fF
C38 a_n29_n430# a_215_n174# 0.13fF
C39 out vdd 0.54fF
C40 a_n29_n330# a_n29_n630# 0.07fF
C41 a_n29_279# a_n29_n330# 0.01fF
C42 a_n29_0# a_n29_679# 0.03fF
C43 a_n29_479# a_n124_86# 0.07fF
C44 a_n29_479# w_n171_117# 0.01fF
C45 a_n29_n330# a_15_n174# 0.14fF
C46 a_n29_n49# vdd 0.01fF
C47 a_n29_n330# out 0.00fF
C48 a_n29_379# a_n124_86# 0.06fF
C49 a_315_n174# a_n29_n49# 0.14fF
C50 a_n29_n730# a_n29_679# 0.01fF
C51 a_n29_379# w_n171_117# 0.01fF
C52 a_n29_n530# a_215_n174# 0.13fF
C53 a_n29_n330# a_n29_n49# 0.01fF
C54 a_515_n174# a_n29_679# 0.13fF
C55 a_n29_n430# a_n29_n730# 0.03fF
C56 a_n29_n430# gnd 1.48fF
C57 a_415_n174# a_215_n174# 0.06fF
C58 a_n29_479# a_n29_379# 0.52fF
C59 a_415_n174# a_n29_779# 0.03fF
C60 a_n29_279# a_115_n174# 0.14fF
C61 a_n29_579# a_n29_679# 0.27fF
C62 a_n29_n630# in 0.08fF
C63 a_215_n174# w_n171_117# 0.00fF
C64 a_415_n174# a_n29_0# 0.01fF
C65 a_n29_n430# a_n29_n230# 0.20fF
C66 a_15_n174# a_115_n174# 0.17fF
C67 w_n171_117# a_n29_779# 0.05fF
C68 a_15_n174# in 0.01fF
C69 a_n29_0# a_n124_86# 0.09fF
C70 a_n29_n530# a_n29_n730# 0.14fF
C71 a_n29_n530# gnd 1.55fF
C72 a_n29_0# w_n171_117# 0.00fF
C73 a_n29_n430# a_n29_n830# 0.01fF
C74 a_n29_479# a_215_n174# 0.13fF
C75 a_n29_479# a_n29_779# 0.01fF
C76 a_115_n174# a_n29_n49# 0.15fF
C77 a_415_n174# a_n29_n730# 0.12fF
C78 a_415_n174# gnd 0.01fF
C79 a_n29_n49# in 0.02fF
C80 a_n29_679# vdd 1.78fF
C81 a_n29_479# a_n29_0# 0.08fF
C82 a_515_n174# a_415_n174# 0.17fF
C83 a_n29_n530# a_n29_n230# 0.09fF
C84 a_n29_379# a_215_n174# 0.13fF
C85 a_n124_86# gnd 1.29fF
C86 a_n29_279# a_15_n174# 0.14fF
C87 a_n29_679# a_315_n174# 0.03fF
C88 a_n29_279# out 0.00fF
C89 a_515_n174# w_n171_117# 0.00fF
C90 a_n29_379# a_n29_779# 0.01fF
C91 a_n29_n530# a_n29_n830# 0.01fF
C92 a_415_n174# a_n29_n230# 0.02fF
C93 a_n29_0# a_n29_379# 0.22fF
C94 a_415_n174# a_n29_579# 0.13fF
C95 a_n29_n430# a_315_n174# 0.03fF
C96 a_n29_n630# a_n29_n49# 0.01fF
C97 a_n29_279# a_n29_n49# 0.01fF
C98 a_n29_n330# a_n29_n430# 0.43fF
C99 a_n124_86# a_n29_n230# 0.08fF
C100 a_415_n174# a_n29_n830# 0.03fF
C101 a_n29_579# a_n124_86# 0.10fF
C102 a_n29_579# w_n171_117# 0.01fF
C103 a_15_n174# a_n29_n49# 0.20fF
C104 a_n29_n49# out 0.32fF
C105 a_n29_0# a_215_n174# 0.01fF
C106 a_n29_479# a_n29_579# 0.58fF
C107 a_415_n174# vdd 0.03fF
C108 a_n29_n530# a_315_n174# 0.13fF
C109 a_n29_0# a_n29_779# 0.01fF
C110 a_n29_n330# a_n29_n530# 0.23fF
C111 a_n124_86# vdd 2.33fF
C112 a_415_n174# a_315_n174# 0.17fF
C113 w_n171_117# vdd 0.07fF
C114 a_415_n174# a_n29_n330# 0.00fF
C115 a_n29_579# a_n29_379# 0.27fF
C116 a_215_n174# gnd 0.01fF
C117 a_n29_n430# a_115_n174# 0.13fF
C118 w_n171_117# a_315_n174# 0.00fF
C119 a_n29_n430# in 0.05fF
C120 a_n29_n330# a_n124_86# 0.03fF
C121 a_n29_479# vdd 1.63fF
C122 a_515_n174# a_n29_779# 0.12fF
C123 a_n29_479# a_315_n174# 0.13fF
C124 a_n29_n230# a_215_n174# 0.03fF
C125 a_n29_279# a_n29_679# 0.03fF
C126 a_n29_579# a_215_n174# 0.03fF
C127 a_n29_379# vdd 1.57fF
C128 a_n29_n430# a_n29_n630# 0.25fF
C129 a_n29_579# a_n29_779# 0.12fF
C130 a_n29_n530# a_115_n174# 0.03fF
C131 a_n29_0# a_n29_n230# 0.01fF
C132 a_n29_n730# gnd 1.79fF
C133 a_n29_n530# in 0.06fF
C134 a_n29_679# out 0.15fF
C135 a_n29_579# a_n29_0# 0.08fF
C136 a_n29_n830# a_n29_779# 0.01fF
C137 a_n29_379# a_315_n174# 0.03fF
C138 a_515_n174# a_n29_n730# 0.13fF
C139 a_n29_n430# a_15_n174# 0.03fF
C140 a_515_n174# gnd 0.00fF
C141 a_415_n174# in 0.00fF
C142 a_n29_679# a_n29_n49# 0.03fF
C143 a_215_n174# vdd 0.03fF
C144 a_115_n174# w_n171_117# 0.00fF
C145 a_n29_n730# a_n29_n230# 0.02fF
C146 a_n29_n230# gnd 0.73fF
C147 a_n124_86# in 0.06fF
C148 a_n29_n430# a_n29_n49# 0.01fF
C149 a_n29_n530# a_n29_n630# 0.55fF
C150 a_n29_779# vdd 3.01fF
C151 a_515_n174# a_n29_579# 0.03fF
C152 a_215_n174# a_315_n174# 0.17fF
C153 a_n29_0# vdd 1.51fF
C154 a_n29_n730# a_n29_n830# 1.30fF
C155 a_n29_n830# gnd 2.09fF
C156 a_n29_479# a_115_n174# 0.03fF
C157 a_n29_n330# a_215_n174# 0.03fF
C158 a_415_n174# a_n29_n630# 0.13fF
C159 a_n29_279# a_415_n174# 0.00fF
C160 a_515_n174# a_n29_n830# 0.15fF
C161 a_n29_0# a_315_n174# 0.01fF
C162 a_n124_86# a_n29_n630# 0.01fF
C163 a_n29_279# a_n124_86# 0.07fF
C164 a_n29_279# w_n171_117# 0.00fF
C165 a_415_n174# out 0.00fF
C166 a_n29_n230# a_n29_n830# 0.01fF
C167 a_n29_n530# a_n29_n49# 0.01fF
C168 a_n29_379# a_115_n174# 0.13fF
C169 a_15_n174# a_n124_86# 0.09fF
C170 a_515_n174# vdd 0.00fF
C171 a_15_n174# w_n171_117# 0.00fF
C172 a_n29_279# a_n29_479# 0.24fF
C173 a_415_n174# a_n29_n49# 0.20fF
C174 w_n171_117# out 0.00fF
C175 a_n29_n730# a_315_n174# 0.03fF
C176 a_315_n174# gnd 0.01fF
C177 a_n29_n330# a_n29_n730# 0.03fF
C178 a_515_n174# a_315_n174# 0.06fF
C179 a_n29_n330# gnd 1.32fF
C180 a_n124_86# a_n29_n49# 0.03fF
C181 w_n171_117# a_n29_n49# 0.00fF
C182 a_n29_479# out 0.00fF
C183 a_n29_579# vdd 1.70fF
C184 a_115_n174# a_215_n174# 0.17fF
C185 a_n29_279# a_n29_379# 0.46fF
C186 a_n29_n230# a_315_n174# 0.03fF
C187 a_n29_479# a_n29_n49# 0.01fF
C188 a_n29_579# a_315_n174# 0.13fF
C189 a_n29_n330# a_n29_n230# 0.33fF
C190 a_n29_0# a_115_n174# 0.04fF
C191 a_15_n174# a_n29_379# 0.03fF
C192 a_n29_379# out 0.00fF
C193 a_n29_n330# a_n29_n830# 0.01fF
C194 a_n29_n630# a_215_n174# 0.03fF
C195 a_n29_279# a_215_n174# 0.03fF
C196 a_n29_379# a_n29_n49# 0.01fF
C197 a_n29_279# a_n29_779# 0.01fF
C198 a_115_n174# gnd 0.01fF
C199 a_15_n174# a_215_n174# 0.06fF
C200 a_315_n174# vdd 0.03fF
C201 gnd in 0.96fF
C202 a_n29_279# a_n29_0# 0.40fF
C203 a_n29_n430# a_n29_n530# 0.49fF
C204 a_415_n174# a_n29_679# 0.12fF
C205 out a_n29_779# 0.27fF
C206 a_n29_0# a_15_n174# 0.14fF
C207 a_115_n174# a_n29_n230# 0.06fF
C208 a_n29_n330# a_315_n174# 0.00fF
C209 a_215_n174# a_n29_n49# 0.14fF
C210 a_n29_0# out 0.00fF
C211 a_n29_n230# in 0.01fF
C212 a_n29_679# w_n171_117# 0.04fF
C213 a_n29_n49# a_n29_779# 0.13fF
C214 a_n29_n730# a_n29_n630# 0.27fF
C215 a_n29_n630# gnd 1.62fF
C216 gnd SUB 3.23fF
C217 in SUB 1.31fF
C218 out SUB 0.62fF
C219 vdd SUB 2.75fF
C220 a_n29_n830# SUB 0.90fF
C221 a_n29_n730# SUB 0.69fF
C222 a_n29_n630# SUB 0.03fF
C223 a_n29_n530# SUB 0.03fF
C224 a_n29_n430# SUB 0.04fF
C225 a_n29_n330# SUB 0.04fF
C226 a_n29_n230# SUB 0.05fF
C227 a_515_n174# SUB 0.30fF
C228 a_415_n174# SUB 0.30fF
C229 a_315_n174# SUB 0.30fF
C230 a_215_n174# SUB 0.30fF
C231 a_115_n174# SUB 0.30fF
C232 a_15_n174# SUB 0.30fF
C233 a_n29_0# SUB 0.04fF
C234 a_n29_279# SUB 0.04fF
C235 a_n29_379# SUB 0.04fF
C236 a_n29_479# SUB 0.02fF
C237 a_n29_n49# SUB 2.12fF
C238 a_n29_579# SUB 0.02fF
C239 a_n29_679# SUB 0.70fF
C240 a_n124_86# SUB 1.55fF
C241 a_n29_779# SUB 0.90fF
C242 w_n171_117# SUB 7.98fF

v1 vdd gnd 1.8
.ends vco


*FD
.subckt fd Clk_In Clk_Out

XM1000 a_79_75# Clk_In VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2088 pd=202 as=1824 ps=170.667
XM1001 GND a_597_66# a_787_62# GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=912 pd=110.667 as=1116 ps=134
XM1002 a_332_67# a_79_75# a_190_75# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=126.737
XM1003 a_463_74# a_332_67# VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2088 pd=217.263 as=1824 ps=170.667
XM1004 a_79_75# Clk_In GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=130 as=912 ps=110.667
XM1005 a_190_75# a_143_127# GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=106.8 as=912 ps=110.667
XM1006 a_143_127# a_597_66# VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2088 pd=202 as=1824 ps=170.667
XM1007 a_597_66# a_79_75# a_463_74# GND sky130_fd_pr__nfet_01v8 w=84 l=15
+  ad=2436 pd=226 as=2436 ps=249.2
XM1008 a_143_127# a_597_66# GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=130 as=912 ps=110.667
XM1009 VDD a_597_66# a_787_62# VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=1824 pd=170.667 as=2232 ps=206
XM1010 Clk_Out a_787_62# GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=130 as=912 ps=110.667
XM1011 a_190_75# a_143_127# VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2088 pd=217.263 as=1824 ps=170.667
XM1012 a_332_67# Clk_In a_190_75# GND sky130_fd_pr__nfet_01v8 w=84 l=15
+  ad=2436 pd=226 as=2436 ps=249.2
XM1013 a_597_66# Clk_In a_463_74# VDD sky130_fd_pr__pfet_01v8 w=42 l=15
+  ad=1218 pd=142 as=1218 ps=126.737
XM1014 Clk_Out a_787_62# VDD VDD sky130_fd_pr__pfet_01v8 w=72 l=15
+  ad=2143 pd=204 as=1824 ps=170.667
XM1015 a_463_74# a_332_67# GND GND sky130_fd_pr__nfet_01v8 w=36 l=15
+  ad=1044 pd=106.8 as=912 ps=110.667
C0 VDD a_143_127# 0.38fF
C1 VDD Clk_Out 0.10fF
C2 a_332_67# a_463_74# 0.12fF
C3 a_332_67# a_190_75# 0.28fF
C4 Clk_Out a_143_127# 0.04fF
C5 VDD a_79_75# 0.37fF
C6 Clk_In a_597_66# 0.17fF
C7 a_79_75# a_143_127# 0.84fF
C8 VDD a_463_74# 0.19fF
C9 VDD a_190_75# 0.22fF
C10 a_463_74# a_143_127# 0.21fF
C11 a_190_75# a_143_127# 0.20fF
C12 VDD a_787_62# 0.21fF
C13 a_463_74# a_79_75# 0.12fF
C14 a_787_62# a_143_127# 0.12fF
C15 a_190_75# a_79_75# 0.29fF
C16 Clk_Out a_787_62# 0.17fF
C17 Clk_In a_332_67# 0.14fF
C18 a_463_74# a_190_75# 0.04fF
C19 a_332_67# a_597_66# 0.02fF
C20 VDD Clk_In 1.10fF
C21 VDD a_597_66# 0.19fF
C22 Clk_In a_143_127# 1.17fF
C23 a_597_66# a_143_127# 0.64fF
C24 Clk_Out a_597_66# 0.01fF
C25 Clk_In a_79_75# 0.60fF
C26 a_597_66# a_79_75# 0.03fF
C27 Clk_In a_463_74# 0.20fF
C28 Clk_In a_190_75# 0.30fF
C29 a_463_74# a_597_66# 0.32fF
C30 VDD a_332_67# 0.15fF
C31 Clk_In a_787_62# 0.01fF
C32 a_332_67# a_143_127# 0.19fF
C33 a_787_62# a_597_66# 0.44fF
C34 a_332_67# a_79_75# 0.16fF
C35 VDD GND 3.76fF
C36 a_787_62# GND 0.47fF
C37 a_597_66# GND 1.33fF
C38 a_463_74# GND 0.36fF
C39 a_332_67# GND 0.44fF
C40 a_190_75# GND 0.38fF
C41 a_79_75# GND 1.06fF
C42 a_143_127# GND 0.99fF 


*c1 7 0 18f
v1 VDD GND 1.8
.ends fd