VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CP
  CLASS CORE ;
  FOREIGN CP ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.670 BY 6.400 ;
  SITE unithddb1 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.120 4.670 20.660 6.260 ;
        RECT 0.120 4.360 8.160 4.670 ;
        RECT 1.960 4.230 8.160 4.360 ;
        RECT 2.300 4.080 8.160 4.230 ;
        RECT 2.410 4.030 8.160 4.080 ;
        RECT 11.580 3.930 20.660 4.670 ;
        RECT 11.580 3.890 19.420 3.930 ;
        RECT 11.580 3.880 12.880 3.890 ;
        RECT 11.580 3.580 12.510 3.880 ;
      LAYER li1 ;
        RECT 0.000 6.070 20.660 6.240 ;
        RECT 2.480 5.850 20.480 6.070 ;
        RECT 13.380 4.200 20.150 4.410 ;
      LAYER mcon ;
        RECT 0.210 6.070 0.380 6.240 ;
        RECT 0.550 6.070 0.720 6.240 ;
        RECT 0.890 6.070 1.060 6.240 ;
        RECT 1.230 6.070 1.400 6.240 ;
        RECT 1.570 6.070 1.740 6.240 ;
        RECT 1.910 6.070 2.080 6.240 ;
        RECT 2.250 6.070 2.420 6.240 ;
        RECT 2.590 6.070 2.760 6.240 ;
        RECT 2.930 6.070 3.100 6.240 ;
        RECT 3.270 6.070 3.440 6.240 ;
        RECT 3.610 6.070 3.780 6.240 ;
        RECT 3.950 6.070 4.120 6.240 ;
        RECT 4.290 6.070 4.460 6.240 ;
        RECT 4.630 6.070 4.800 6.240 ;
        RECT 4.970 6.070 5.140 6.240 ;
        RECT 5.310 6.070 5.480 6.240 ;
        RECT 5.650 6.070 5.820 6.240 ;
        RECT 5.990 6.070 6.160 6.240 ;
        RECT 6.330 6.070 6.500 6.240 ;
        RECT 6.670 6.070 6.840 6.240 ;
        RECT 7.010 6.070 7.180 6.240 ;
        RECT 7.350 6.070 7.520 6.240 ;
        RECT 7.690 6.070 7.860 6.240 ;
        RECT 8.030 6.070 8.200 6.240 ;
        RECT 8.370 6.070 8.540 6.240 ;
        RECT 8.710 6.070 8.880 6.240 ;
        RECT 9.050 6.070 9.220 6.240 ;
        RECT 9.390 6.070 9.560 6.240 ;
        RECT 9.730 6.070 9.900 6.240 ;
        RECT 10.070 6.070 10.240 6.240 ;
        RECT 10.410 6.070 10.580 6.240 ;
        RECT 10.750 6.070 10.920 6.240 ;
        RECT 11.090 6.070 11.260 6.240 ;
        RECT 11.430 6.070 11.600 6.240 ;
        RECT 11.770 6.070 11.940 6.240 ;
        RECT 12.110 6.070 12.280 6.240 ;
        RECT 12.450 6.070 12.620 6.240 ;
        RECT 12.790 6.070 12.960 6.240 ;
        RECT 13.130 6.070 13.300 6.240 ;
        RECT 13.470 6.070 13.640 6.240 ;
        RECT 13.810 6.070 13.980 6.240 ;
        RECT 14.150 6.070 14.320 6.240 ;
        RECT 14.490 6.070 14.660 6.240 ;
        RECT 14.830 6.070 15.000 6.240 ;
        RECT 15.170 6.070 15.340 6.240 ;
        RECT 15.510 6.070 15.680 6.240 ;
        RECT 15.850 6.070 16.020 6.240 ;
        RECT 16.190 6.070 16.360 6.240 ;
        RECT 16.530 6.070 16.700 6.240 ;
        RECT 16.870 6.070 17.040 6.240 ;
        RECT 17.210 6.070 17.380 6.240 ;
        RECT 17.550 6.070 17.720 6.240 ;
        RECT 17.890 6.070 18.060 6.240 ;
        RECT 18.230 6.070 18.400 6.240 ;
        RECT 18.570 6.070 18.740 6.240 ;
        RECT 18.910 6.070 19.080 6.240 ;
        RECT 19.250 6.070 19.420 6.240 ;
        RECT 19.590 6.070 19.760 6.240 ;
        RECT 19.930 6.070 20.100 6.240 ;
        RECT 20.270 6.070 20.440 6.240 ;
        RECT 18.820 4.220 18.990 4.390 ;
        RECT 19.250 4.220 19.420 4.390 ;
      LAYER met1 ;
        RECT 0.000 5.920 20.660 6.400 ;
        RECT 18.760 4.460 19.460 5.920 ;
        RECT 18.760 4.160 19.480 4.460 ;
    END
    PORT
      LAYER nwell ;
        RECT 0.600 1.170 3.150 1.680 ;
        RECT 0.600 0.320 3.900 1.170 ;
        RECT 10.550 1.150 11.390 1.600 ;
        RECT 10.550 0.310 12.410 1.150 ;
      LAYER li1 ;
        RECT 3.220 0.320 3.900 0.730 ;
        RECT 11.600 0.320 12.410 0.820 ;
        RECT 0.000 0.150 20.670 0.320 ;
      LAYER mcon ;
        RECT 0.210 0.150 0.380 0.320 ;
        RECT 0.550 0.150 0.720 0.320 ;
        RECT 0.890 0.150 1.060 0.320 ;
        RECT 1.230 0.150 1.400 0.320 ;
        RECT 1.570 0.150 1.740 0.320 ;
        RECT 1.910 0.150 2.080 0.320 ;
        RECT 2.250 0.150 2.420 0.320 ;
        RECT 2.590 0.150 2.760 0.320 ;
        RECT 2.930 0.150 3.100 0.320 ;
        RECT 3.270 0.150 3.440 0.320 ;
        RECT 3.610 0.150 3.780 0.320 ;
        RECT 3.950 0.150 4.120 0.320 ;
        RECT 4.290 0.150 4.460 0.320 ;
        RECT 4.630 0.150 4.800 0.320 ;
        RECT 4.970 0.150 5.140 0.320 ;
        RECT 5.310 0.150 5.480 0.320 ;
        RECT 5.650 0.150 5.820 0.320 ;
        RECT 5.990 0.150 6.160 0.320 ;
        RECT 6.330 0.150 6.500 0.320 ;
        RECT 6.670 0.150 6.840 0.320 ;
        RECT 7.010 0.150 7.180 0.320 ;
        RECT 7.350 0.150 7.520 0.320 ;
        RECT 7.690 0.150 7.860 0.320 ;
        RECT 8.030 0.150 8.200 0.320 ;
        RECT 8.370 0.150 8.540 0.320 ;
        RECT 8.710 0.150 8.880 0.320 ;
        RECT 9.050 0.150 9.220 0.320 ;
        RECT 9.390 0.150 9.560 0.320 ;
        RECT 9.730 0.150 9.900 0.320 ;
        RECT 10.070 0.150 10.240 0.320 ;
        RECT 10.410 0.150 10.580 0.320 ;
        RECT 10.750 0.150 10.920 0.320 ;
        RECT 11.090 0.150 11.260 0.320 ;
        RECT 11.430 0.150 11.600 0.320 ;
        RECT 11.770 0.150 11.940 0.320 ;
        RECT 12.110 0.150 12.280 0.320 ;
        RECT 12.450 0.150 12.620 0.320 ;
        RECT 12.790 0.150 12.960 0.320 ;
        RECT 13.130 0.150 13.300 0.320 ;
        RECT 13.470 0.150 13.640 0.320 ;
        RECT 13.810 0.150 13.980 0.320 ;
        RECT 14.150 0.150 14.320 0.320 ;
        RECT 14.490 0.150 14.660 0.320 ;
        RECT 14.830 0.150 15.000 0.320 ;
        RECT 15.170 0.150 15.340 0.320 ;
        RECT 15.510 0.150 15.680 0.320 ;
        RECT 15.850 0.150 16.020 0.320 ;
        RECT 16.190 0.150 16.360 0.320 ;
        RECT 16.530 0.150 16.700 0.320 ;
        RECT 16.870 0.150 17.040 0.320 ;
        RECT 17.210 0.150 17.380 0.320 ;
        RECT 17.550 0.150 17.720 0.320 ;
        RECT 17.890 0.150 18.060 0.320 ;
        RECT 18.230 0.150 18.400 0.320 ;
        RECT 18.570 0.150 18.740 0.320 ;
        RECT 18.910 0.150 19.080 0.320 ;
        RECT 19.250 0.150 19.420 0.320 ;
        RECT 19.590 0.150 19.760 0.320 ;
        RECT 19.930 0.150 20.100 0.320 ;
      LAYER met1 ;
        RECT 0.000 0.000 20.670 0.480 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.300 3.270 6.370 3.550 ;
        RECT 8.600 3.270 9.020 3.520 ;
        RECT 0.010 3.100 10.410 3.270 ;
        RECT 11.140 3.100 20.660 3.270 ;
        RECT 0.930 2.040 1.120 3.100 ;
        RECT 2.170 2.040 2.360 3.100 ;
        RECT 4.010 2.730 9.250 3.100 ;
        RECT 12.080 2.820 19.570 3.100 ;
        RECT 4.010 2.720 9.420 2.730 ;
        RECT 3.880 2.550 9.420 2.720 ;
        RECT 4.620 2.540 9.420 2.550 ;
      LAYER mcon ;
        RECT 0.210 3.100 0.380 3.270 ;
        RECT 0.550 3.100 0.720 3.270 ;
        RECT 0.890 3.100 1.060 3.270 ;
        RECT 1.230 3.100 1.400 3.270 ;
        RECT 1.570 3.100 1.740 3.270 ;
        RECT 1.910 3.100 2.080 3.270 ;
        RECT 2.250 3.100 2.420 3.270 ;
        RECT 2.590 3.100 2.760 3.270 ;
        RECT 2.930 3.100 3.100 3.270 ;
        RECT 3.270 3.100 3.440 3.270 ;
        RECT 3.610 3.100 3.780 3.270 ;
        RECT 3.950 3.100 4.120 3.270 ;
        RECT 4.290 3.100 4.460 3.270 ;
        RECT 4.630 3.100 4.800 3.270 ;
        RECT 4.970 3.100 5.140 3.270 ;
        RECT 5.310 3.100 5.480 3.270 ;
        RECT 5.650 3.100 5.820 3.270 ;
        RECT 5.990 3.100 6.160 3.270 ;
        RECT 6.330 3.100 6.500 3.270 ;
        RECT 6.670 3.100 6.840 3.270 ;
        RECT 7.010 3.100 7.180 3.270 ;
        RECT 7.350 3.100 7.520 3.270 ;
        RECT 7.690 3.100 7.860 3.270 ;
        RECT 8.030 3.100 8.200 3.270 ;
        RECT 8.370 3.100 8.540 3.270 ;
        RECT 8.710 3.100 8.880 3.270 ;
        RECT 9.050 3.100 9.220 3.270 ;
        RECT 9.390 3.100 9.560 3.270 ;
        RECT 9.730 3.100 9.900 3.270 ;
        RECT 10.070 3.100 10.240 3.270 ;
        RECT 11.430 3.100 11.600 3.270 ;
        RECT 11.770 3.100 11.940 3.270 ;
        RECT 12.110 3.100 12.280 3.270 ;
        RECT 12.450 3.100 12.620 3.270 ;
        RECT 12.790 3.100 12.960 3.270 ;
        RECT 13.130 3.100 13.300 3.270 ;
        RECT 13.470 3.100 13.640 3.270 ;
        RECT 13.810 3.100 13.980 3.270 ;
        RECT 14.150 3.100 14.320 3.270 ;
        RECT 14.490 3.100 14.660 3.270 ;
        RECT 14.830 3.100 15.000 3.270 ;
        RECT 15.170 3.100 15.340 3.270 ;
        RECT 15.510 3.100 15.680 3.270 ;
        RECT 15.850 3.100 16.020 3.270 ;
        RECT 16.190 3.100 16.360 3.270 ;
        RECT 16.530 3.100 16.700 3.270 ;
        RECT 16.870 3.100 17.040 3.270 ;
        RECT 17.210 3.100 17.380 3.270 ;
        RECT 17.550 3.100 17.720 3.270 ;
        RECT 17.890 3.100 18.060 3.270 ;
        RECT 18.230 3.100 18.400 3.270 ;
        RECT 18.570 3.100 18.740 3.270 ;
        RECT 18.910 3.100 19.080 3.270 ;
        RECT 19.250 3.100 19.420 3.270 ;
        RECT 19.590 3.100 19.760 3.270 ;
        RECT 19.930 3.100 20.100 3.270 ;
      LAYER met1 ;
        RECT 0.010 2.960 20.660 3.440 ;
    END
  END GND
  PIN Up
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.225000 ;
    PORT
      LAYER li1 ;
        RECT 10.100 2.490 10.270 2.820 ;
        RECT 1.940 1.660 2.270 1.830 ;
      LAYER mcon ;
        RECT 10.100 2.570 10.270 2.740 ;
        RECT 2.020 1.660 2.190 1.830 ;
      LAYER met1 ;
        RECT 10.020 2.490 10.340 2.810 ;
        RECT 1.940 1.580 2.260 1.900 ;
      LAYER via ;
        RECT 10.050 2.520 10.310 2.780 ;
        RECT 1.970 1.610 2.230 1.870 ;
      LAYER met2 ;
        RECT 9.470 2.490 10.340 2.810 ;
        RECT 1.760 1.610 2.260 1.900 ;
        RECT 1.760 1.100 2.090 1.610 ;
        RECT 9.470 1.100 9.840 2.490 ;
        RECT 1.760 1.090 9.840 1.100 ;
        RECT 0.010 0.730 9.840 1.090 ;
    END
  END Up
  PIN Down
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.972000 ;
    PORT
      LAYER li1 ;
        RECT 2.040 4.030 2.210 4.360 ;
        RECT 0.700 1.660 1.030 1.830 ;
      LAYER mcon ;
        RECT 2.040 4.110 2.210 4.280 ;
        RECT 0.780 1.660 0.950 1.830 ;
      LAYER met1 ;
        RECT 1.960 4.030 2.280 4.350 ;
        RECT 0.710 1.580 1.030 1.900 ;
      LAYER via ;
        RECT 1.990 4.060 2.250 4.320 ;
        RECT 0.740 1.610 1.000 1.870 ;
      LAYER met2 ;
        RECT 1.840 4.330 2.280 4.350 ;
        RECT 0.600 4.030 2.280 4.330 ;
        RECT 0.600 3.970 2.270 4.030 ;
        RECT 0.600 2.720 0.920 3.970 ;
        RECT 0.010 2.410 0.920 2.720 ;
        RECT 0.600 1.900 0.920 2.410 ;
        RECT 0.600 1.580 1.030 1.900 ;
    END
  END Down
  PIN Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.277200 ;
    PORT
      LAYER li1 ;
        RECT 11.850 3.870 20.660 4.020 ;
        RECT 10.610 3.490 20.660 3.870 ;
        RECT 10.610 3.480 11.960 3.490 ;
        RECT 10.610 2.730 10.960 3.480 ;
        RECT 10.540 2.560 10.960 2.730 ;
    END
  END Out
  PIN ENb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.700000 ;
    PORT
      LAYER li1 ;
        RECT 0.510 4.810 0.960 5.050 ;
    END
  END ENb
  OBS
      LAYER li1 ;
        RECT 1.720 5.390 20.480 5.580 ;
        RECT 8.370 5.340 8.750 5.390 ;
        RECT 9.630 5.340 10.010 5.390 ;
        RECT 11.870 5.340 12.250 5.390 ;
        RECT 1.220 4.900 2.160 5.090 ;
        RECT 2.480 4.900 20.480 5.090 ;
        RECT 8.370 4.850 8.750 4.900 ;
        RECT 9.630 4.850 10.010 4.900 ;
        RECT 2.480 4.350 9.020 4.520 ;
        RECT 11.870 4.500 12.250 4.900 ;
        RECT 7.990 3.760 8.240 4.350 ;
        RECT 8.430 4.300 9.020 4.350 ;
        RECT 11.850 4.310 12.270 4.500 ;
        RECT 8.480 4.250 9.020 4.300 ;
        RECT 8.550 4.190 9.020 4.250 ;
        RECT 8.600 3.830 9.020 4.190 ;
        RECT 11.220 4.080 11.550 4.250 ;
        RECT 7.950 3.590 8.280 3.760 ;
        RECT 1.410 2.500 1.670 2.760 ;
        RECT 0.930 0.690 1.120 1.450 ;
        RECT 1.410 0.730 1.600 2.500 ;
        RECT 2.650 1.740 2.840 2.400 ;
        RECT 3.370 2.060 4.320 2.250 ;
        RECT 10.540 2.220 10.960 2.250 ;
        RECT 9.990 2.170 10.960 2.220 ;
        RECT 4.620 1.980 10.960 2.170 ;
        RECT 2.170 0.700 2.360 1.460 ;
        RECT 2.650 1.380 4.310 1.740 ;
        RECT 4.620 1.500 11.150 1.690 ;
        RECT 2.650 0.740 2.840 1.380 ;
        RECT 10.170 1.100 10.420 1.500 ;
        RECT 10.600 1.460 11.150 1.500 ;
        RECT 10.670 1.420 11.150 1.460 ;
        RECT 10.720 1.370 11.150 1.420 ;
        RECT 10.730 1.170 11.150 1.370 ;
        RECT 10.130 0.930 10.460 1.100 ;
        RECT 10.730 0.690 11.150 0.900 ;
      LAYER mcon ;
        RECT 12.810 5.400 12.980 5.570 ;
        RECT 13.150 5.400 13.320 5.570 ;
        RECT 11.300 4.080 11.470 4.250 ;
        RECT 1.460 2.540 1.630 2.710 ;
        RECT 0.940 1.110 1.110 1.280 ;
        RECT 0.940 0.770 1.110 0.940 ;
        RECT 2.180 1.120 2.350 1.290 ;
        RECT 2.180 0.780 2.350 0.950 ;
        RECT 10.860 0.720 11.030 0.890 ;
      LAYER met1 ;
        RECT 12.750 5.340 13.430 5.630 ;
        RECT 11.220 4.020 11.540 4.320 ;
        RECT 1.380 2.460 1.700 2.780 ;
        RECT 12.680 1.540 13.470 2.290 ;
        RECT 0.900 0.990 1.150 1.340 ;
        RECT 2.140 0.990 2.390 1.350 ;
        RECT 12.680 0.990 13.160 1.540 ;
        RECT 0.900 0.690 13.160 0.990 ;
      LAYER via ;
        RECT 12.930 5.340 13.190 5.600 ;
        RECT 11.250 4.030 11.510 4.290 ;
        RECT 1.410 2.490 1.670 2.750 ;
        RECT 12.810 1.740 13.350 2.100 ;
      LAYER met2 ;
        RECT 8.700 4.000 11.540 4.320 ;
        RECT 8.700 3.000 9.170 4.000 ;
        RECT 1.380 2.600 9.170 3.000 ;
        RECT 1.380 2.460 1.700 2.600 ;
        RECT 12.780 1.710 13.390 5.630 ;
  END
END CP
MACRO VCO_new
  CLASS BLOCK ;
  FOREIGN VCO_new ;
  ORIGIN 1.740 9.100 ;
  SIZE 8.950 BY 17.540 ;
  PIN in
    ANTENNAGATEAREA 6.000000 ;
    PORT
      LAYER li1 ;
        RECT -1.740 -1.710 -1.330 -1.540 ;
    END
  END in
  PIN vdd
    ANTENNADIFFAREA 12.818000 ;
    PORT
      LAYER li1 ;
        RECT -0.630 8.190 6.700 8.440 ;
        RECT -0.630 7.580 -0.460 8.190 ;
        RECT -0.630 7.410 4.710 7.580 ;
        RECT -0.630 7.020 -0.460 7.410 ;
        RECT -1.590 6.850 -0.460 7.020 ;
        RECT -1.470 1.350 -1.300 6.850 ;
        RECT -0.630 6.580 -0.460 6.850 ;
        RECT -0.630 6.410 4.710 6.580 ;
        RECT -0.630 5.580 -0.460 6.410 ;
        RECT -0.630 5.410 4.710 5.580 ;
        RECT -0.630 4.580 -0.460 5.410 ;
        RECT -0.630 4.410 4.710 4.580 ;
        RECT -0.630 3.580 -0.460 4.410 ;
        RECT -0.630 3.410 4.710 3.580 ;
        RECT -0.630 2.580 -0.460 3.410 ;
        RECT -0.630 2.410 4.710 2.580 ;
        RECT -0.630 1.580 -0.460 2.410 ;
        RECT 5.770 1.590 5.940 8.190 ;
        RECT -0.630 1.410 4.600 1.580 ;
      LAYER mcon ;
        RECT -0.550 8.230 -0.380 8.400 ;
        RECT -0.180 8.230 -0.010 8.400 ;
        RECT 0.260 8.230 0.430 8.400 ;
        RECT 0.710 8.230 0.880 8.400 ;
        RECT 1.150 8.230 1.320 8.400 ;
        RECT 1.590 8.230 1.760 8.400 ;
        RECT 2.040 8.230 2.210 8.400 ;
        RECT 2.480 8.230 2.650 8.400 ;
        RECT 2.920 8.230 3.090 8.400 ;
        RECT 3.360 8.230 3.530 8.400 ;
        RECT 3.810 8.230 3.980 8.400 ;
        RECT 4.250 8.230 4.420 8.400 ;
        RECT 4.690 8.230 4.860 8.400 ;
        RECT 5.140 8.230 5.310 8.400 ;
        RECT 5.580 8.230 5.750 8.400 ;
        RECT 6.020 8.230 6.190 8.400 ;
        RECT 6.470 8.230 6.640 8.400 ;
        RECT -0.630 7.810 -0.460 7.980 ;
        RECT -0.630 7.450 -0.460 7.620 ;
        RECT -0.630 7.040 -0.460 7.210 ;
        RECT -1.390 6.850 -1.220 7.020 ;
        RECT -0.990 6.850 -0.820 7.020 ;
        RECT -0.630 6.620 -0.460 6.790 ;
        RECT -0.630 6.190 -0.460 6.360 ;
        RECT -0.630 5.770 -0.460 5.940 ;
        RECT -0.630 5.340 -0.460 5.510 ;
        RECT -0.630 4.920 -0.460 5.090 ;
        RECT -0.630 4.490 -0.460 4.660 ;
        RECT -0.630 4.070 -0.460 4.240 ;
        RECT -0.630 3.640 -0.460 3.810 ;
        RECT -0.630 3.220 -0.460 3.390 ;
        RECT -0.630 2.790 -0.460 2.960 ;
        RECT -0.630 2.370 -0.460 2.540 ;
        RECT -0.630 1.930 -0.460 2.100 ;
      LAYER met1 ;
        RECT -0.670 8.190 6.700 8.440 ;
        RECT -0.670 7.060 -0.420 8.190 ;
        RECT -1.470 6.810 -0.420 7.060 ;
        RECT -0.670 1.350 -0.420 6.810 ;
    END
  END vdd
  PIN gnd
    ANTENNADIFFAREA 11.913199 ;
    PORT
      LAYER li1 ;
        RECT -1.470 -7.510 -1.300 -2.010 ;
        RECT -0.670 -2.510 -0.420 -2.430 ;
        RECT -0.670 -2.630 4.710 -2.510 ;
        RECT -0.630 -2.680 4.710 -2.630 ;
        RECT -0.630 -3.510 -0.460 -2.680 ;
        RECT -0.630 -3.680 4.710 -3.510 ;
        RECT -0.630 -4.510 -0.460 -3.680 ;
        RECT -0.630 -4.680 4.710 -4.510 ;
        RECT -0.630 -5.510 -0.460 -4.680 ;
        RECT -0.630 -5.680 4.710 -5.510 ;
        RECT -0.630 -6.510 -0.460 -5.680 ;
        RECT -0.630 -6.680 4.710 -6.510 ;
        RECT -0.630 -7.510 -0.460 -6.680 ;
        RECT -1.590 -7.680 4.710 -7.510 ;
        RECT -0.630 -8.510 -0.460 -7.680 ;
        RECT 5.770 -8.510 5.940 -2.250 ;
        RECT -0.630 -8.680 5.940 -8.510 ;
        RECT -0.630 -8.850 -0.460 -8.680 ;
        RECT -0.210 -8.850 -0.040 -8.680 ;
        RECT 0.240 -8.850 0.410 -8.680 ;
        RECT 0.630 -8.850 0.800 -8.680 ;
        RECT 1.020 -8.850 1.190 -8.680 ;
        RECT 1.470 -8.850 1.640 -8.680 ;
        RECT 1.920 -8.850 2.090 -8.680 ;
        RECT 2.370 -8.850 2.540 -8.680 ;
        RECT 2.820 -8.850 2.990 -8.680 ;
        RECT 3.270 -8.850 3.440 -8.680 ;
        RECT 3.710 -8.850 3.880 -8.680 ;
        RECT 4.160 -8.850 4.330 -8.680 ;
        RECT 4.500 -8.850 4.670 -8.680 ;
        RECT -0.630 -9.100 6.760 -8.850 ;
      LAYER mcon ;
        RECT -0.630 -2.660 -0.460 -2.490 ;
        RECT -0.630 -3.120 -0.460 -2.950 ;
        RECT -0.630 -3.580 -0.460 -3.410 ;
        RECT -0.630 -4.050 -0.460 -3.880 ;
        RECT -0.630 -4.970 -0.460 -4.800 ;
        RECT -0.630 -5.440 -0.460 -5.270 ;
        RECT -0.630 -5.900 -0.460 -5.730 ;
        RECT -0.630 -6.360 -0.460 -6.190 ;
        RECT -0.630 -6.830 -0.460 -6.660 ;
        RECT -0.630 -7.290 -0.460 -7.120 ;
        RECT -1.390 -7.680 -1.220 -7.510 ;
        RECT -0.990 -7.680 -0.820 -7.510 ;
        RECT -0.630 -7.750 -0.460 -7.580 ;
        RECT -0.630 -8.220 -0.460 -8.050 ;
        RECT -0.550 -9.070 -0.380 -8.900 ;
        RECT -0.060 -9.070 0.110 -8.900 ;
        RECT 0.550 -9.070 0.720 -8.900 ;
        RECT 1.170 -9.070 1.340 -8.900 ;
        RECT 1.780 -9.070 1.950 -8.900 ;
        RECT 2.400 -9.070 2.570 -8.900 ;
        RECT 3.010 -9.070 3.180 -8.900 ;
        RECT 3.630 -9.070 3.800 -8.900 ;
        RECT 4.240 -9.070 4.410 -8.900 ;
        RECT 4.860 -9.070 5.030 -8.900 ;
        RECT 5.470 -9.070 5.640 -8.900 ;
        RECT 6.090 -9.070 6.260 -8.900 ;
        RECT 6.530 -9.060 6.700 -8.890 ;
      LAYER met1 ;
        RECT -0.670 -7.470 -0.420 -2.430 ;
        RECT -1.470 -7.720 -0.420 -7.470 ;
        RECT -0.670 -8.850 -0.420 -7.720 ;
        RECT -0.670 -9.100 6.760 -8.850 ;
    END
  END gnd
  PIN out
    ANTENNADIFFAREA 1.531200 ;
    PORT
      LAYER li1 ;
        RECT 6.210 1.840 6.380 5.790 ;
        RECT 6.150 1.670 7.030 1.840 ;
        RECT 6.210 1.590 6.380 1.670 ;
        RECT 6.860 -0.240 7.030 1.670 ;
        RECT 6.860 -0.410 7.210 -0.240 ;
        RECT 6.210 -2.330 6.380 -2.250 ;
        RECT 6.860 -2.330 7.030 -0.410 ;
        RECT 6.150 -2.500 7.030 -2.330 ;
        RECT 6.210 -3.330 6.380 -2.500 ;
    END
  END out
  OBS
      LAYER nwell ;
        RECT -0.470 6.530 6.620 8.260 ;
        RECT -1.710 1.170 6.620 6.530 ;
        RECT -0.470 -0.180 6.620 1.170 ;
      LAYER li1 ;
        RECT -0.290 7.850 5.560 8.020 ;
        RECT -0.290 6.850 5.050 7.020 ;
        RECT -1.030 -7.010 -0.860 6.350 ;
        RECT -0.290 5.850 4.710 6.020 ;
        RECT -0.290 4.850 4.710 5.020 ;
        RECT -0.290 3.850 4.710 4.020 ;
        RECT -0.290 2.850 4.710 3.020 ;
        RECT -0.290 1.850 4.710 2.020 ;
        RECT 4.880 1.420 5.050 6.850 ;
        RECT 4.770 1.250 5.050 1.420 ;
        RECT 5.390 1.420 5.560 7.850 ;
        RECT 5.390 1.250 5.940 1.420 ;
        RECT -0.230 0.000 -0.060 1.080 ;
        RECT 0.210 -0.250 0.380 1.080 ;
        RECT 0.770 0.000 0.940 1.080 ;
        RECT 1.210 -0.250 1.380 1.080 ;
        RECT 1.770 0.000 1.940 1.080 ;
        RECT 2.210 -0.250 2.380 1.080 ;
        RECT 2.770 0.000 2.940 1.080 ;
        RECT 3.210 -0.250 3.380 1.080 ;
        RECT 3.770 0.000 3.940 1.080 ;
        RECT 4.210 -0.250 4.380 1.080 ;
        RECT 4.770 0.000 4.940 1.250 ;
        RECT 5.210 -0.250 5.380 1.080 ;
        RECT 5.770 0.000 5.940 1.250 ;
        RECT 6.210 -0.240 6.380 1.080 ;
        RECT -0.290 -0.420 0.040 -0.250 ;
        RECT 0.210 -0.420 1.040 -0.250 ;
        RECT 1.210 -0.420 2.040 -0.250 ;
        RECT 2.210 -0.420 3.040 -0.250 ;
        RECT 3.210 -0.420 4.040 -0.250 ;
        RECT 4.210 -0.420 5.040 -0.250 ;
        RECT 5.210 -0.420 6.040 -0.250 ;
        RECT 6.210 -0.410 6.690 -0.240 ;
        RECT -0.230 -2.070 -0.060 -0.660 ;
        RECT 0.210 -1.740 0.380 -0.420 ;
        RECT 0.770 -1.740 0.940 -0.660 ;
        RECT 1.210 -1.740 1.380 -0.420 ;
        RECT 1.770 -1.740 1.940 -0.660 ;
        RECT 2.210 -1.740 2.380 -0.420 ;
        RECT 2.770 -1.740 2.940 -0.660 ;
        RECT 3.210 -1.740 3.380 -0.420 ;
        RECT 3.770 -1.740 3.940 -0.660 ;
        RECT 4.210 -1.740 4.380 -0.420 ;
        RECT 4.770 -1.910 4.940 -0.660 ;
        RECT 5.210 -1.740 5.380 -0.420 ;
        RECT 5.770 -1.910 5.940 -0.660 ;
        RECT 6.210 -1.740 6.380 -0.410 ;
        RECT -0.290 -2.240 4.600 -2.070 ;
        RECT 4.770 -2.080 5.050 -1.910 ;
        RECT -0.290 -3.240 4.710 -3.070 ;
        RECT -0.290 -4.240 4.710 -4.070 ;
        RECT -0.290 -5.240 4.710 -5.070 ;
        RECT -0.290 -6.240 4.710 -6.070 ;
        RECT 4.880 -7.070 5.050 -2.080 ;
        RECT -0.290 -7.240 5.050 -7.070 ;
        RECT 5.220 -2.080 5.940 -1.910 ;
        RECT 5.220 -8.070 5.390 -2.080 ;
        RECT -0.290 -8.240 5.390 -8.070 ;
      LAYER mcon ;
        RECT 3.850 5.850 4.020 6.020 ;
        RECT 2.760 4.850 2.930 5.020 ;
        RECT 1.660 3.850 1.830 4.020 ;
        RECT 0.900 2.850 1.070 3.020 ;
        RECT -0.130 1.850 0.040 2.020 ;
        RECT -0.230 0.910 -0.060 1.080 ;
        RECT 0.770 0.910 0.940 1.080 ;
        RECT 1.770 0.910 1.940 1.080 ;
        RECT 2.770 0.910 2.940 1.080 ;
        RECT 3.770 0.910 3.940 1.080 ;
        RECT -0.290 -0.420 -0.120 -0.250 ;
        RECT 6.360 -0.410 6.530 -0.240 ;
        RECT 0.770 -3.240 0.940 -3.070 ;
        RECT 1.790 -4.240 1.960 -4.070 ;
        RECT 2.780 -5.240 2.950 -5.070 ;
        RECT 3.780 -6.240 3.950 -6.070 ;
      LAYER met1 ;
        RECT 3.710 5.790 4.110 6.080 ;
        RECT 1.570 3.790 2.000 4.080 ;
        RECT 0.710 2.790 1.150 3.080 ;
        RECT -0.280 1.790 0.110 2.080 ;
        RECT -0.280 0.830 -0.010 1.790 ;
        RECT 0.710 0.830 1.000 2.790 ;
        RECT 1.710 0.830 2.000 3.790 ;
        RECT 2.710 0.830 3.000 5.080 ;
        RECT 3.710 0.830 4.000 5.790 ;
        RECT -0.470 -0.490 6.620 -0.180 ;
        RECT 0.710 -3.300 1.000 -1.490 ;
        RECT 1.710 -4.300 2.000 -1.490 ;
        RECT 2.710 -5.300 3.000 -1.490 ;
        RECT 3.710 -6.300 4.000 -1.490 ;
  END
END VCO_new
MACRO PFD
  CLASS CORE ;
  FOREIGN PFD ;
  ORIGIN 0.000 0.000 ;
  SIZE 7.670 BY 6.400 ;
  SITE unithddb1 ;
  PIN Clk_Ref
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.879000 ;
    ANTENNADIFFAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 2.420 5.520 3.520 5.710 ;
        RECT 2.420 5.210 2.650 5.520 ;
        RECT 0.040 1.740 0.310 3.510 ;
        RECT 0.040 1.450 2.100 1.740 ;
    END
  END Clk_Ref
  PIN Up
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.427200 ;
    PORT
      LAYER li1 ;
        RECT 6.270 4.780 6.560 5.780 ;
        RECT 6.390 4.040 6.560 4.780 ;
        RECT 6.260 3.560 6.560 4.040 ;
    END
  END Up
  PIN Down
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.427200 ;
    PORT
      LAYER li1 ;
        RECT 6.520 1.930 6.810 2.930 ;
        RECT 6.640 1.190 6.810 1.930 ;
        RECT 6.510 0.710 6.810 1.190 ;
    END
  END Down
  PIN Clk2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.879000 ;
    ANTENNADIFFAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 0.900 2.060 1.230 2.230 ;
        RECT 4.700 1.850 4.890 2.720 ;
        RECT 4.390 1.620 4.890 1.850 ;
      LAYER mcon ;
        RECT 0.980 2.060 1.150 2.230 ;
      LAYER met1 ;
        RECT 0.710 2.010 1.210 2.290 ;
    END
  END Clk2
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 4.340 3.290 5.010 4.100 ;
        RECT 5.780 3.360 6.000 3.880 ;
        RECT 5.560 3.290 6.230 3.360 ;
        RECT 4.340 3.120 7.670 3.290 ;
        RECT 0.780 2.760 0.990 2.780 ;
        RECT 0.700 2.590 1.060 2.760 ;
        RECT 0.780 2.510 0.990 2.590 ;
        RECT 1.730 0.920 1.910 1.280 ;
        RECT 6.030 0.700 6.250 1.030 ;
      LAYER mcon ;
        RECT 4.940 3.120 5.110 3.290 ;
        RECT 5.280 3.120 5.450 3.290 ;
        RECT 5.620 3.120 5.790 3.290 ;
        RECT 5.960 3.120 6.130 3.290 ;
        RECT 6.300 3.120 6.470 3.290 ;
        RECT 6.640 3.120 6.810 3.290 ;
        RECT 0.800 2.590 0.970 2.760 ;
        RECT 1.740 1.010 1.910 1.180 ;
        RECT 6.070 0.780 6.240 0.950 ;
      LAYER met1 ;
        RECT 0.000 2.960 7.670 3.440 ;
        RECT 0.740 2.530 1.040 2.960 ;
        RECT 2.280 1.240 2.520 2.960 ;
        RECT 1.680 0.950 2.520 1.240 ;
        RECT 5.600 1.010 5.870 2.960 ;
        RECT 5.600 0.720 6.270 1.010 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.890 5.350 7.670 6.400 ;
        RECT 1.370 4.790 7.670 5.350 ;
        RECT 5.050 4.600 7.670 4.790 ;
      LAYER li1 ;
        RECT 0.000 6.050 7.670 6.220 ;
        RECT 1.650 5.720 2.070 6.050 ;
        RECT 1.510 5.510 2.220 5.720 ;
        RECT 5.770 5.080 6.000 6.050 ;
      LAYER mcon ;
        RECT 0.800 6.050 0.970 6.220 ;
        RECT 1.140 6.050 1.310 6.220 ;
        RECT 1.480 6.050 1.650 6.220 ;
        RECT 1.820 6.050 1.990 6.220 ;
        RECT 2.160 6.050 2.330 6.220 ;
        RECT 2.500 6.050 2.670 6.220 ;
        RECT 2.840 6.050 3.010 6.220 ;
        RECT 3.180 6.050 3.350 6.220 ;
        RECT 3.520 6.050 3.690 6.220 ;
        RECT 3.860 6.050 4.030 6.220 ;
        RECT 4.200 6.050 4.370 6.220 ;
        RECT 4.540 6.050 4.710 6.220 ;
        RECT 4.880 6.050 5.050 6.220 ;
        RECT 5.220 6.050 5.390 6.220 ;
        RECT 5.560 6.050 5.730 6.220 ;
        RECT 5.900 6.050 6.070 6.220 ;
        RECT 6.240 6.050 6.410 6.220 ;
        RECT 6.580 6.050 6.750 6.220 ;
      LAYER met1 ;
        RECT 0.000 5.920 7.670 6.400 ;
    END
    PORT
      LAYER nwell ;
        RECT 6.770 3.070 7.670 3.080 ;
        RECT 4.430 2.950 7.670 3.070 ;
        RECT 3.970 1.570 7.670 2.950 ;
        RECT 3.970 0.310 5.140 1.570 ;
      LAYER li1 ;
        RECT 6.020 2.540 6.250 2.930 ;
        RECT 7.040 2.660 7.450 2.830 ;
        RECT 6.020 2.250 6.330 2.540 ;
        RECT 7.100 2.370 7.400 2.660 ;
        RECT 6.020 2.230 6.250 2.250 ;
        RECT 7.040 2.200 7.450 2.370 ;
        RECT 7.100 1.930 7.400 2.200 ;
        RECT 7.040 1.760 7.450 1.930 ;
        RECT 4.690 0.310 4.900 1.420 ;
        RECT 0.000 0.140 7.670 0.310 ;
      LAYER mcon ;
        RECT 6.160 2.310 6.330 2.480 ;
        RECT 7.140 2.180 7.350 2.390 ;
        RECT 0.800 0.140 0.970 0.310 ;
        RECT 1.140 0.140 1.310 0.310 ;
        RECT 1.480 0.140 1.650 0.310 ;
        RECT 1.820 0.140 1.990 0.310 ;
        RECT 2.160 0.140 2.330 0.310 ;
        RECT 2.500 0.140 2.670 0.310 ;
        RECT 2.840 0.140 3.010 0.310 ;
        RECT 3.180 0.140 3.350 0.310 ;
        RECT 3.520 0.140 3.690 0.310 ;
        RECT 3.860 0.140 4.030 0.310 ;
        RECT 4.200 0.140 4.370 0.310 ;
        RECT 4.540 0.140 4.710 0.310 ;
        RECT 4.880 0.140 5.050 0.310 ;
        RECT 5.220 0.140 5.390 0.310 ;
        RECT 5.560 0.140 5.730 0.310 ;
        RECT 5.900 0.140 6.070 0.310 ;
        RECT 6.240 0.140 6.410 0.310 ;
        RECT 6.580 0.140 6.750 0.310 ;
      LAYER met1 ;
        RECT 6.100 2.250 7.410 2.540 ;
        RECT 6.560 2.070 7.410 2.250 ;
        RECT 6.560 0.480 6.860 2.070 ;
        RECT 0.000 0.000 7.670 0.480 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT 1.550 4.880 2.240 5.240 ;
        RECT 0.370 4.630 2.240 4.880 ;
        RECT 2.840 5.040 3.550 5.230 ;
        RECT 0.370 3.950 0.640 4.630 ;
        RECT 2.840 4.570 3.280 5.040 ;
        RECT 5.260 4.910 5.480 5.780 ;
        RECT 5.260 4.740 6.100 4.910 ;
        RECT 5.900 4.610 6.100 4.740 ;
        RECT 2.840 4.450 5.710 4.570 ;
        RECT 0.870 4.400 5.710 4.450 ;
        RECT 0.870 4.190 3.290 4.400 ;
        RECT 5.900 4.270 6.130 4.610 ;
        RECT 5.900 4.230 6.090 4.270 ;
        RECT 5.250 4.060 6.090 4.230 ;
        RECT 0.370 3.710 3.100 3.950 ;
        RECT 5.250 3.680 5.470 4.060 ;
        RECT 2.860 0.860 3.050 3.320 ;
        RECT 3.340 2.510 3.530 3.320 ;
        RECT 4.220 2.620 4.410 2.750 ;
        RECT 3.950 2.510 4.410 2.620 ;
        RECT 3.340 2.260 4.410 2.510 ;
        RECT 3.340 2.200 3.640 2.260 ;
        RECT 3.340 1.090 3.600 2.200 ;
        RECT 3.950 2.180 4.410 2.260 ;
        RECT 4.220 2.070 4.410 2.180 ;
        RECT 5.510 2.060 5.730 2.930 ;
        RECT 5.510 1.890 6.350 2.060 ;
        RECT 6.160 1.760 6.350 1.890 ;
        RECT 5.140 1.550 5.960 1.720 ;
        RECT 6.160 1.470 6.380 1.760 ;
        RECT 3.340 0.860 3.530 1.090 ;
        RECT 3.960 0.750 4.420 1.440 ;
        RECT 6.150 1.420 6.380 1.470 ;
        RECT 6.150 1.380 6.330 1.420 ;
        RECT 5.500 1.210 6.330 1.380 ;
        RECT 5.500 0.830 5.720 1.210 ;
      LAYER mcon ;
        RECT 2.870 1.240 3.040 1.410 ;
        RECT 3.430 2.230 3.600 2.400 ;
        RECT 5.200 1.550 5.370 1.720 ;
        RECT 4.090 1.000 4.260 1.170 ;
      LAYER met1 ;
        RECT 3.340 2.140 3.690 2.490 ;
        RECT 5.130 1.470 5.450 1.790 ;
        RECT 2.810 1.230 3.790 1.470 ;
        RECT 2.810 1.180 4.320 1.230 ;
        RECT 3.560 0.940 4.320 1.180 ;
      LAYER via ;
        RECT 3.370 2.170 3.660 2.460 ;
        RECT 5.160 1.500 5.420 1.760 ;
      LAYER met2 ;
        RECT 3.340 2.460 3.690 2.490 ;
        RECT 3.340 2.190 5.400 2.460 ;
        RECT 3.340 2.140 3.690 2.190 ;
        RECT 5.140 1.790 5.400 2.190 ;
        RECT 5.130 1.470 5.450 1.790 ;
  END
END PFD
MACRO FD
  CLASS CORE ;
  FOREIGN FD ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.350 BY 3.200 ;
  SITE unithddb1 ;
  PIN Clk_Out
    ANTENNADIFFAREA 0.318700 ;
    PORT
      LAYER li1 ;
        RECT 8.910 2.550 9.090 2.590 ;
        RECT 8.910 1.810 9.200 2.550 ;
        RECT 8.950 1.640 9.200 1.810 ;
        RECT 9.030 0.980 9.200 1.640 ;
        RECT 8.900 0.620 9.200 0.980 ;
    END
  END Clk_Out
  PIN GND
    ANTENNADIFFAREA 1.261200 ;
    PORT
      LAYER li1 ;
        RECT 0.410 0.320 0.580 1.110 ;
        RECT 1.520 0.320 1.690 1.110 ;
        RECT 4.250 0.320 4.420 1.100 ;
        RECT 6.910 0.320 7.080 1.110 ;
        RECT 8.420 0.320 8.640 0.910 ;
        RECT 0.000 0.150 9.350 0.320 ;
      LAYER mcon ;
        RECT 0.160 0.150 0.330 0.320 ;
        RECT 1.000 0.150 1.170 0.320 ;
        RECT 1.800 0.150 1.970 0.320 ;
        RECT 3.150 0.150 3.320 0.320 ;
        RECT 4.070 0.150 4.240 0.320 ;
        RECT 5.130 0.150 5.300 0.320 ;
        RECT 5.970 0.150 6.140 0.320 ;
        RECT 7.150 0.150 7.320 0.320 ;
        RECT 7.990 0.150 8.160 0.320 ;
        RECT 8.830 0.150 9.000 0.320 ;
      LAYER met1 ;
        RECT 0.000 0.000 9.350 0.480 ;
    END
  END GND
  PIN Clk_In
    ANTENNAGATEAREA 0.351000 ;
    PORT
      LAYER li1 ;
        RECT 6.490 2.160 6.660 2.500 ;
        RECT 0.000 1.310 0.660 1.480 ;
        RECT 2.370 0.740 2.700 0.920 ;
      LAYER mcon ;
        RECT 6.490 2.240 6.660 2.410 ;
        RECT 0.410 1.310 0.580 1.480 ;
        RECT 2.450 0.750 2.620 0.920 ;
      LAYER met1 ;
        RECT 0.350 2.180 1.570 2.500 ;
        RECT 6.440 2.490 6.720 2.500 ;
        RECT 0.350 1.270 0.640 2.180 ;
        RECT 1.320 2.070 1.570 2.180 ;
        RECT 6.430 2.070 6.720 2.490 ;
        RECT 1.320 1.820 6.720 2.070 ;
        RECT 0.360 0.980 0.640 1.270 ;
        RECT 0.360 0.690 2.710 0.980 ;
    END
  END Clk_In
  PIN VDD
    ANTENNADIFFAREA 1.829700 ;
    PORT
      LAYER nwell ;
        RECT 0.000 1.850 9.320 3.200 ;
        RECT 0.000 1.490 2.370 1.850 ;
        RECT 3.960 1.840 9.320 1.850 ;
        RECT 3.960 1.490 5.100 1.840 ;
        RECT 6.670 1.600 9.320 1.840 ;
        RECT 6.670 1.550 7.860 1.600 ;
        RECT 6.790 1.480 7.860 1.550 ;
      LAYER li1 ;
        RECT 0.000 2.830 9.320 3.020 ;
        RECT 0.410 1.730 0.580 2.830 ;
        RECT 1.520 1.730 1.690 2.830 ;
        RECT 4.250 1.720 4.420 2.830 ;
        RECT 6.910 1.730 7.080 2.830 ;
        RECT 8.410 2.220 8.640 2.830 ;
      LAYER mcon ;
        RECT 0.550 2.830 0.740 3.020 ;
        RECT 1.370 2.830 1.560 3.020 ;
        RECT 2.820 2.830 3.010 3.020 ;
        RECT 3.600 2.830 3.790 3.020 ;
        RECT 4.540 2.830 4.730 3.020 ;
        RECT 5.620 2.830 5.810 3.020 ;
        RECT 6.820 2.830 7.010 3.020 ;
        RECT 7.680 2.830 7.870 3.020 ;
        RECT 8.540 2.830 8.730 3.020 ;
      LAYER met1 ;
        RECT 0.000 2.720 9.320 3.200 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT 0.850 1.560 1.020 2.450 ;
        RECT 1.960 1.570 2.130 2.450 ;
        RECT 2.440 2.220 2.610 2.550 ;
        RECT 2.940 1.930 3.110 2.460 ;
        RECT 2.390 1.630 3.110 1.930 ;
        RECT 2.390 1.570 2.640 1.630 ;
        RECT 0.850 1.260 1.150 1.560 ;
        RECT 1.430 1.310 1.770 1.480 ;
        RECT 1.960 1.270 2.640 1.570 ;
        RECT 0.850 0.750 1.020 1.260 ;
        RECT 1.960 0.750 2.130 1.270 ;
        RECT 2.940 0.830 3.110 1.630 ;
        RECT 3.380 1.900 3.550 2.460 ;
        RECT 3.380 1.630 4.080 1.900 ;
        RECT 3.380 0.830 3.550 1.630 ;
        RECT 3.910 1.540 4.080 1.630 ;
        RECT 4.690 1.560 4.860 2.440 ;
        RECT 5.590 1.910 5.760 2.450 ;
        RECT 5.090 1.620 5.760 1.910 ;
        RECT 5.090 1.560 5.370 1.620 ;
        RECT 3.910 1.520 4.120 1.540 ;
        RECT 3.910 1.470 4.460 1.520 ;
        RECT 3.910 1.300 4.500 1.470 ;
        RECT 3.910 1.270 4.460 1.300 ;
        RECT 4.690 1.270 5.370 1.560 ;
        RECT 4.690 0.740 4.860 1.270 ;
        RECT 5.090 0.710 5.420 0.880 ;
        RECT 5.590 0.820 5.760 1.620 ;
        RECT 6.030 1.880 6.200 2.450 ;
        RECT 6.030 1.630 6.570 1.880 ;
        RECT 6.030 0.820 6.200 1.630 ;
        RECT 6.380 1.520 6.570 1.630 ;
        RECT 7.350 1.560 7.520 2.450 ;
        RECT 7.900 2.010 8.120 2.590 ;
        RECT 7.900 1.840 8.740 2.010 ;
        RECT 8.550 1.640 8.740 1.840 ;
        RECT 6.790 1.520 7.120 1.530 ;
        RECT 6.380 1.480 7.120 1.520 ;
        RECT 6.380 1.310 7.160 1.480 ;
        RECT 6.380 1.280 7.120 1.310 ;
        RECT 6.380 1.010 6.570 1.280 ;
        RECT 7.350 1.260 7.690 1.560 ;
        RECT 8.010 1.420 8.350 1.590 ;
        RECT 8.550 1.350 8.770 1.640 ;
        RECT 8.540 1.300 8.770 1.350 ;
        RECT 6.380 0.700 6.660 1.010 ;
        RECT 7.350 0.750 7.520 1.260 ;
        RECT 8.540 1.250 8.720 1.300 ;
        RECT 7.890 1.080 8.720 1.250 ;
        RECT 7.890 0.620 8.110 1.080 ;
      LAYER mcon ;
        RECT 2.440 2.290 2.610 2.470 ;
        RECT 0.910 1.320 1.080 1.490 ;
        RECT 1.520 1.310 1.690 1.480 ;
        RECT 5.170 0.710 5.340 0.880 ;
        RECT 7.440 1.320 7.610 1.490 ;
        RECT 8.100 1.420 8.270 1.590 ;
        RECT 6.460 0.770 6.630 0.940 ;
      LAYER met1 ;
        RECT 2.370 2.220 2.690 2.540 ;
        RECT 0.830 1.240 1.180 1.590 ;
        RECT 1.460 1.260 7.690 1.540 ;
        RECT 8.040 1.370 8.350 1.650 ;
        RECT 8.070 1.000 8.340 1.370 ;
        RECT 5.080 0.630 5.410 0.960 ;
        RECT 6.400 0.730 8.340 1.000 ;
        RECT 6.400 0.710 6.720 0.730 ;
        RECT 6.410 0.700 6.720 0.710 ;
      LAYER via ;
        RECT 2.400 2.250 2.660 2.510 ;
        RECT 0.880 1.290 1.140 1.550 ;
        RECT 5.110 0.660 5.380 0.930 ;
      LAYER met2 ;
        RECT 0.850 1.590 1.180 1.660 ;
        RECT 0.830 1.570 1.180 1.590 ;
        RECT 2.370 1.570 2.690 2.510 ;
        RECT 0.830 1.280 5.400 1.570 ;
        RECT 0.830 1.240 1.180 1.280 ;
        RECT 5.070 0.930 5.400 1.280 ;
        RECT 5.070 0.870 5.410 0.930 ;
        RECT 5.080 0.630 5.410 0.870 ;
  END
END FD
MACRO MUX
  CLASS CORE ;
  FOREIGN MUX ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.080 BY 2.970 ;
  SITE unithddb1 ;
  PIN SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.324000 ;
    PORT
      LAYER li1 ;
        RECT 2.760 2.630 3.090 2.800 ;
        RECT 0.760 0.370 1.090 0.540 ;
        RECT 1.630 0.350 1.960 0.560 ;
      LAYER mcon ;
        RECT 2.840 2.630 3.010 2.800 ;
        RECT 0.840 0.370 1.010 0.540 ;
        RECT 1.710 0.370 1.880 0.540 ;
      LAYER met1 ;
        RECT 2.760 2.550 3.080 2.870 ;
        RECT 1.630 0.600 1.950 0.610 ;
        RECT 0.000 0.300 1.950 0.600 ;
        RECT 1.630 0.290 1.950 0.300 ;
      LAYER via ;
        RECT 2.790 2.580 3.050 2.840 ;
        RECT 1.660 0.320 1.920 0.580 ;
      LAYER met2 ;
        RECT 2.760 2.830 3.080 2.870 ;
        RECT 2.230 2.580 3.080 2.830 ;
        RECT 1.630 0.600 1.950 0.610 ;
        RECT 2.230 0.600 2.480 2.580 ;
        RECT 2.760 2.550 3.080 2.580 ;
        RECT 1.630 0.300 2.480 0.600 ;
        RECT 1.630 0.290 1.950 0.300 ;
    END
  END SEL
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.313200 ;
    PORT
      LAYER li1 ;
        RECT 2.610 0.740 2.780 2.340 ;
      LAYER mcon ;
        RECT 2.610 2.120 2.780 2.290 ;
      LAYER met1 ;
        RECT 0.000 2.060 2.840 2.350 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.313200 ;
    PORT
      LAYER li1 ;
        RECT 1.480 1.490 1.650 2.340 ;
        RECT 1.330 1.220 1.650 1.490 ;
        RECT 1.480 0.740 1.650 1.220 ;
      LAYER mcon ;
        RECT 1.350 1.260 1.520 1.430 ;
      LAYER met1 ;
        RECT 0.000 1.200 1.580 1.500 ;
    END
  END B
  PIN Out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.626400 ;
    PORT
      LAYER li1 ;
        RECT 1.920 0.740 2.090 2.340 ;
        RECT 3.050 2.320 3.220 2.340 ;
        RECT 3.050 2.090 3.340 2.320 ;
        RECT 3.050 0.740 3.220 2.090 ;
      LAYER mcon ;
        RECT 1.920 1.280 2.090 1.450 ;
        RECT 3.140 2.120 3.310 2.290 ;
      LAYER met1 ;
        RECT 3.080 2.060 3.900 2.350 ;
        RECT 3.630 1.880 3.900 2.060 ;
        RECT 3.630 1.510 4.080 1.880 ;
        RECT 1.860 1.460 4.080 1.510 ;
        RECT 1.860 1.220 3.920 1.460 ;
    END
  END Out
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 0.120 2.520 1.710 2.970 ;
        RECT 0.120 1.440 3.460 2.520 ;
      LAYER li1 ;
        RECT 0.420 1.620 0.590 2.930 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.420 0.200 0.590 1.100 ;
        RECT 0.300 0.000 0.710 0.200 ;
    END
  END GND
  OBS
      LAYER li1 ;
        RECT 0.860 2.610 2.440 2.820 ;
        RECT 0.860 0.740 1.030 2.610 ;
        RECT 2.270 0.570 2.440 2.610 ;
        RECT 2.270 0.360 3.090 0.570 ;
  END
END MUX
END LIBRARY

