magic
tech sky130A
timestamp 1633597695
<< error_s >>
rect -1706 1538 -1691 1544
rect -1655 1538 -1640 1544
rect -1551 1525 -1536 1531
rect -1285 1526 -1270 1532
rect -1012 1525 -997 1531
rect -901 1525 -886 1531
rect -1706 1496 -1691 1502
rect -1655 1496 -1640 1502
rect -1551 1483 -1536 1489
rect -1285 1484 -1270 1490
rect -1012 1483 -997 1489
rect -901 1483 -886 1489
rect -1512 1376 -1507 1400
rect -1488 1359 -1483 1376
rect -1448 1359 -1447 1397
rect -2225 1201 -2224 1205
rect -2201 1184 -2200 1201
rect -2165 1184 -2160 1205
rect -1132 1201 -1131 1205
rect -1108 1184 -1107 1201
rect -1072 1184 -1067 1205
rect -2786 1071 -2771 1077
rect -2675 1071 -2660 1077
rect -2402 1070 -2387 1076
rect -2136 1071 -2121 1077
rect -1693 1071 -1678 1077
rect -1582 1071 -1567 1077
rect -1309 1070 -1294 1076
rect -1043 1071 -1028 1077
rect -2032 1058 -2017 1064
rect -1981 1058 -1966 1064
rect -939 1058 -924 1064
rect -888 1058 -873 1064
rect -2786 1029 -2771 1035
rect -2675 1029 -2660 1035
rect -2402 1028 -2387 1034
rect -2136 1029 -2121 1035
rect -1693 1029 -1678 1035
rect -1582 1029 -1567 1035
rect -1309 1028 -1294 1034
rect -1043 1029 -1028 1035
rect -2032 1016 -2017 1022
rect -1981 1016 -1966 1022
rect -939 1016 -924 1022
rect -888 1016 -873 1022
rect -2799 898 -2784 904
rect -2748 898 -2733 904
rect -1706 898 -1691 904
rect -1655 898 -1640 904
rect -2644 885 -2629 891
rect -2378 886 -2363 892
rect -2105 885 -2090 891
rect -1994 885 -1979 891
rect -1551 885 -1536 891
rect -1285 886 -1270 892
rect -1012 885 -997 891
rect -901 885 -886 891
rect -2799 856 -2784 862
rect -2748 856 -2733 862
rect -1706 856 -1691 862
rect -1655 856 -1640 862
rect -2644 843 -2629 849
rect -2378 844 -2363 850
rect -2105 843 -2090 849
rect -1994 843 -1979 849
rect -1551 843 -1536 849
rect -1285 844 -1270 850
rect -1012 843 -997 849
rect -901 843 -886 849
rect -1608 800 -1568 812
rect -2605 736 -2600 760
rect -2581 719 -2576 736
rect -2541 719 -2540 757
rect -1512 736 -1507 760
rect -1488 719 -1483 736
rect -1448 719 -1447 757
rect -2755 605 -2753 622
rect -2736 605 -2722 622
rect -2721 605 -2719 622
rect -2702 605 -2700 622
rect -2687 605 -2685 622
rect -2668 605 -2666 622
rect -2653 605 -2640 622
rect -2634 605 -2632 622
rect -2619 605 -2617 622
rect -2600 605 -2598 622
rect -2585 605 -2583 622
rect -2570 605 -2558 622
rect -2551 605 -2549 622
rect -2532 605 -2530 622
rect -2517 605 -2515 622
rect -2498 605 -2496 622
rect -2488 605 -2476 622
rect -2464 605 -2462 622
rect -2449 605 -2447 622
rect -2430 605 -2428 622
rect -2415 605 -2413 622
rect -2406 605 -2394 622
rect -2381 605 -2379 622
rect -2362 605 -2360 622
rect -2347 605 -2345 622
rect -2328 605 -2326 622
rect -2313 605 -2311 622
rect -2294 605 -2292 622
rect -2279 605 -2277 622
rect -2260 605 -2258 622
rect -2245 605 -2243 622
rect -2226 605 -2224 622
rect -2211 605 -2209 622
rect -2192 605 -2190 622
rect -2047 607 -2045 624
rect -2028 607 -2026 624
rect -2013 607 -2011 624
rect -1994 607 -1992 624
rect -1979 607 -1977 624
rect -1960 607 -1958 624
rect -1945 607 -1943 624
rect -1926 607 -1924 624
rect -1911 607 -1909 624
rect -1892 607 -1890 624
rect -1877 607 -1875 624
rect -1858 607 -1856 624
rect -1843 607 -1841 624
rect -1824 607 -1822 624
rect -1809 607 -1807 624
rect -1790 607 -1788 624
rect -1775 607 -1773 624
rect -1756 607 -1754 624
rect -1741 607 -1739 624
rect -1722 607 -1720 624
rect -1707 607 -1705 624
rect -1688 607 -1686 624
rect -1673 607 -1671 624
rect -1654 607 -1652 624
rect -1639 607 -1637 624
rect -1620 607 -1618 624
rect -1605 607 -1603 624
rect -1586 607 -1584 624
rect -1571 607 -1569 624
rect -1552 607 -1550 624
rect -1537 607 -1535 624
rect -1518 607 -1516 624
rect -1503 607 -1501 624
rect -1484 607 -1482 624
rect -1469 607 -1467 624
rect -1450 607 -1448 624
rect -1435 607 -1433 624
rect -1416 607 -1414 624
rect -1401 607 -1399 624
rect -1382 607 -1380 624
rect -1367 607 -1365 624
rect -1348 607 -1346 624
rect -1333 607 -1331 624
rect -1314 607 -1312 624
rect -1299 607 -1297 624
rect -1280 607 -1278 624
rect -1265 607 -1263 624
rect -1246 607 -1244 624
rect -1231 607 -1229 624
rect -1212 607 -1210 624
rect -1197 607 -1195 624
rect -1178 607 -1176 624
rect -1163 607 -1161 624
rect -1144 607 -1142 624
rect -1129 607 -1127 624
rect -1110 607 -1108 624
rect -1095 607 -1093 624
rect -1076 607 -1074 624
rect -1061 607 -1059 624
rect -1042 607 -1040 624
rect -1027 607 -1025 624
rect -1008 607 -1006 624
rect -993 607 -991 624
rect -974 607 -972 624
rect -959 607 -957 624
rect -940 607 -938 624
rect -925 607 -923 624
rect -906 607 -904 624
rect -891 607 -889 624
rect -872 607 -870 624
rect -857 607 -855 624
rect -838 607 -836 624
rect -823 607 -821 624
rect -804 607 -802 624
rect -789 607 -787 624
rect -770 607 -768 624
rect -755 607 -753 624
rect -736 607 -734 624
rect -721 607 -719 624
rect -702 607 -700 624
rect -687 607 -685 624
rect -668 607 -666 624
rect -653 607 -651 624
rect -634 607 -632 624
rect -619 607 -617 624
rect -600 607 -598 624
rect -585 607 -583 624
rect -566 607 -564 624
rect -551 607 -549 624
rect -532 607 -530 624
rect -517 607 -515 624
rect -498 607 -496 624
rect -483 607 -481 624
rect -464 607 -462 624
rect -449 607 -447 624
rect -430 607 -428 624
rect -415 607 -413 624
rect -396 607 -394 624
rect -381 607 -379 624
rect -362 607 -360 624
rect -347 607 -345 624
rect -328 607 -326 624
rect -313 607 -311 624
rect -294 607 -292 624
rect -279 607 -277 624
rect -260 607 -258 624
rect -245 607 -243 624
rect -226 607 -224 624
rect -211 607 -209 624
rect -192 607 -190 624
rect -177 607 -175 624
rect -158 607 -156 624
rect -143 607 -141 624
rect -124 607 -122 624
rect -109 607 -107 624
rect -90 607 -88 624
rect -75 607 -73 624
rect -56 607 -54 624
rect -787 540 -785 557
rect -768 540 -766 557
rect -2272 478 -2263 481
rect -2071 460 -1956 461
rect -744 422 -732 439
rect -662 422 -650 439
rect -580 422 -568 439
rect -498 422 -486 439
rect -416 422 -404 439
rect -334 422 -322 439
rect -252 422 -240 439
rect -170 422 -158 439
rect -2296 404 -2281 410
rect -2296 362 -2281 368
rect -1938 332 -1926 349
rect -1856 332 -1844 349
rect -1774 332 -1762 349
rect -1692 332 -1680 349
rect -1610 332 -1598 349
rect -1528 332 -1516 349
rect -2341 312 -2339 329
rect -2322 312 -2320 329
rect -2307 312 -2305 329
rect -2288 312 -2286 329
rect -2273 312 -2271 329
rect -2254 312 -2252 329
rect -2239 312 -2237 329
rect -2220 312 -2218 329
rect -2205 312 -2203 329
rect -2186 312 -2184 329
rect -2047 310 -2045 327
rect -2028 310 -2026 327
rect -2013 310 -2011 327
rect -1994 310 -1992 327
rect -1979 310 -1977 327
rect -1960 310 -1958 327
rect -1945 310 -1943 327
rect -1926 310 -1924 327
rect -1911 310 -1909 327
rect -1892 310 -1890 327
rect -1877 310 -1875 327
rect -1858 310 -1856 327
rect -1843 310 -1841 327
rect -1824 310 -1822 327
rect -1809 310 -1807 327
rect -1790 310 -1788 327
rect -1775 310 -1773 327
rect -1756 310 -1754 327
rect -1741 310 -1739 327
rect -1722 310 -1720 327
rect -1707 310 -1705 327
rect -1688 310 -1686 327
rect -1673 310 -1671 327
rect -1654 310 -1652 327
rect -1639 310 -1637 327
rect -1620 310 -1618 327
rect -1605 310 -1603 327
rect -1586 310 -1584 327
rect -1571 310 -1569 327
rect -1552 310 -1550 327
rect -1537 310 -1535 327
rect -1518 310 -1516 327
rect -1503 310 -1501 327
rect -1484 310 -1482 327
rect -1469 310 -1467 327
rect -1450 310 -1448 327
rect -1435 310 -1433 327
rect -1416 310 -1414 327
rect -1401 310 -1399 327
rect -1382 310 -1380 327
rect -1367 310 -1365 327
rect -1348 310 -1346 327
rect -1333 310 -1331 327
rect -1314 310 -1312 327
rect -1299 310 -1297 327
rect -1280 310 -1278 327
rect -1265 310 -1263 327
rect -1246 310 -1244 327
rect -1231 310 -1229 327
rect -1212 310 -1210 327
rect -1197 310 -1195 327
rect -1178 310 -1176 327
rect -1163 310 -1161 327
rect -1144 310 -1142 327
rect -1129 310 -1127 327
rect -1110 310 -1108 327
rect -1095 310 -1093 327
rect -1076 310 -1074 327
rect -925 310 -923 327
rect -906 310 -904 327
rect -891 310 -889 327
rect -872 310 -870 327
rect -857 310 -855 327
rect -838 310 -836 327
rect -823 310 -821 327
rect -804 310 -802 327
rect -789 310 -787 327
rect -770 310 -768 327
rect -755 310 -753 327
rect -736 310 -734 327
rect -721 310 -719 327
rect -702 310 -700 327
rect -687 310 -685 327
rect -668 310 -666 327
rect -653 310 -651 327
rect -634 310 -632 327
rect -619 310 -617 327
rect -600 310 -598 327
rect -585 310 -583 327
rect -566 310 -564 327
rect -551 310 -549 327
rect -532 310 -530 327
rect -517 310 -515 327
rect -498 310 -496 327
rect -483 310 -481 327
rect -464 310 -462 327
rect -449 310 -447 327
rect -430 310 -428 327
rect -415 310 -413 327
rect -396 310 -394 327
rect -381 310 -379 327
rect -362 310 -360 327
rect -347 310 -345 327
rect -328 310 -326 327
rect -313 310 -311 327
rect -294 310 -292 327
rect -279 310 -277 327
rect -260 310 -258 327
rect -245 310 -243 327
rect -226 310 -224 327
rect -211 310 -209 327
rect -192 310 -190 327
rect -177 310 -175 327
rect -158 310 -156 327
rect -143 310 -141 327
rect -124 310 -122 327
rect -109 310 -107 327
rect -90 310 -88 327
rect -2786 284 -2780 299
rect -2744 284 -2738 299
rect -860 287 -848 304
rect -778 287 -766 304
rect -696 287 -684 304
rect -614 287 -602 304
rect -532 287 -520 304
rect -450 287 -438 304
rect -372 287 -360 304
rect -290 287 -278 304
rect -208 287 -196 304
rect -2146 266 -2134 283
rect -2030 240 -2020 274
rect -1964 240 -1949 246
rect -1840 240 -1825 246
rect -2146 220 -2134 237
rect -1996 204 -1986 240
rect -1964 198 -1949 204
rect -1840 198 -1825 204
rect -2247 193 -2238 196
rect -2146 176 -2134 193
rect -2005 166 -1988 169
rect -1881 166 -1864 170
rect -2651 128 -2636 134
rect -2271 119 -2256 125
rect -2187 122 -2186 136
rect -2199 105 -2186 119
rect -1989 111 -1972 113
rect -1865 112 -1848 114
rect -1989 92 -1972 94
rect -1865 93 -1848 95
rect -2651 86 -2636 92
rect -2271 77 -2256 83
rect -1752 50 -1740 67
rect -915 61 -903 78
rect -2755 14 -2753 31
rect -2736 14 -2734 31
rect -2721 14 -2719 31
rect -2702 14 -2700 31
rect -2687 14 -2685 31
rect -2668 14 -2666 31
rect -2653 14 -2651 31
rect -2634 14 -2632 31
rect -2619 14 -2617 31
rect -2600 14 -2598 31
rect -2585 14 -2583 31
rect -2566 14 -2564 31
rect -2551 14 -2549 31
rect -2532 14 -2530 31
rect -2517 14 -2515 31
rect -2498 14 -2496 31
rect -2483 14 -2481 31
rect -2464 14 -2462 31
rect -2449 14 -2447 31
rect -2430 14 -2428 31
rect -2415 14 -2413 31
rect -2396 14 -2394 31
rect -2381 14 -2379 31
rect -2362 14 -2360 31
rect -2347 14 -2345 31
rect -2328 14 -2326 31
rect -2313 14 -2311 31
rect -2294 14 -2292 31
rect -2279 14 -2277 31
rect -2260 14 -2258 31
rect -2245 14 -2243 31
rect -2226 14 -2224 31
rect -2211 14 -2209 31
rect -2192 14 -2190 31
rect -2047 15 -2045 32
rect -2028 15 -2026 32
rect -2013 15 -2011 32
rect -1994 15 -1992 32
rect -1979 15 -1977 32
rect -1960 15 -1958 32
rect -1945 15 -1943 32
rect -1926 15 -1924 32
rect -1911 15 -1909 32
rect -1892 15 -1890 32
rect -1877 15 -1875 32
rect -1858 15 -1856 32
rect -1843 15 -1841 32
rect -1824 15 -1822 32
rect -1809 15 -1807 32
rect -1790 15 -1788 32
rect -1775 15 -1773 32
rect -1756 15 -1754 32
rect -1741 15 -1739 32
rect -1722 15 -1720 32
rect -1707 15 -1705 32
rect -1688 15 -1686 32
rect -1673 15 -1671 32
rect -1654 15 -1652 32
rect -1639 15 -1637 32
rect -1620 15 -1618 32
rect -1605 15 -1603 32
rect -1586 15 -1584 32
rect -1571 15 -1569 32
rect -1552 15 -1550 32
rect -1537 15 -1535 32
rect -1518 15 -1516 32
rect -1503 15 -1501 32
rect -1484 15 -1482 32
rect -1469 15 -1467 32
rect -1450 15 -1448 32
rect -1435 15 -1433 32
rect -1416 15 -1414 32
rect -1401 15 -1399 32
rect -1382 15 -1380 32
rect -1367 15 -1365 32
rect -1348 15 -1346 32
rect -1333 15 -1331 32
rect -1314 15 -1312 32
rect -1299 15 -1297 32
rect -1280 15 -1278 32
rect -1265 15 -1263 32
rect -1246 15 -1244 32
rect -1231 15 -1229 32
rect -1212 15 -1210 32
rect -1197 15 -1195 32
rect -1178 15 -1176 32
rect -1163 15 -1161 32
rect -1144 15 -1142 32
rect -1129 15 -1127 32
rect -1110 15 -1108 32
rect -1095 15 -1093 32
rect -1076 15 -1074 32
rect -1061 15 -1059 32
rect -1042 15 -1040 32
rect -1027 15 -1025 32
rect -1008 15 -1006 32
rect -993 15 -991 32
rect -974 15 -972 32
rect -959 15 -957 32
rect -940 15 -938 32
rect -925 15 -923 32
rect -906 15 -904 32
rect -891 15 -889 32
rect -872 15 -870 32
rect -857 15 -855 32
rect -838 15 -836 32
rect -823 15 -821 32
rect -804 15 -802 32
rect -789 15 -787 32
rect -770 15 -768 32
rect -755 15 -753 32
rect -736 15 -734 32
rect -721 15 -719 32
rect -702 15 -700 32
rect -687 15 -685 32
rect -668 15 -666 32
rect -653 15 -651 32
rect -634 15 -632 32
rect -619 15 -617 32
rect -600 15 -598 32
rect -585 15 -583 32
rect -566 15 -564 32
rect -551 15 -549 32
rect -532 15 -530 32
rect -517 15 -515 32
rect -498 15 -496 32
rect -483 15 -481 32
rect -464 15 -462 32
rect -449 15 -447 32
rect -430 15 -428 32
rect -415 15 -413 32
rect -396 15 -394 32
rect -381 15 -379 32
rect -362 15 -360 32
rect -347 15 -345 32
rect -328 15 -326 32
rect -313 15 -311 32
rect -294 15 -292 32
rect -279 15 -277 32
rect -260 15 -258 32
rect -245 15 -243 32
rect -226 15 -224 32
rect -211 15 -209 32
rect -192 15 -190 32
rect -177 15 -175 32
rect -158 15 -156 32
rect -143 15 -141 32
rect -124 15 -122 32
rect -109 15 -107 32
rect -90 15 -88 32
<< nwell >>
rect -1964 800 -1695 801
rect -2079 785 -1695 800
rect -2101 753 -1695 785
rect -2101 639 -822 753
rect -2127 593 -822 639
rect -2127 461 -1968 593
rect -2103 168 -2020 308
rect -2104 31 -1956 168
<< locali >>
rect -58 1595 -47 1612
rect -30 1595 -5 1612
rect 12 1595 32 1612
rect -839 1568 -729 1585
rect -58 1576 -38 1595
rect -58 1570 -57 1576
rect -3051 1448 -3021 1462
rect -3051 1418 -2826 1448
rect -3051 1404 -3021 1418
rect -2850 1243 -2826 1418
rect -1808 1444 -1725 1461
rect -848 1452 -784 1469
rect -1808 1341 -1791 1444
rect -1874 1322 -1791 1341
rect -1757 1262 -1735 1317
rect -1939 1243 -1735 1262
rect -801 1111 -784 1452
rect -2894 1091 -2833 1108
rect -1945 1091 -1740 1108
rect -853 1094 -784 1111
rect -2894 826 -2877 1091
rect -1933 973 -1915 987
rect -1757 973 -1739 990
rect -1933 969 -1739 973
rect -1933 952 -1853 969
rect -1836 952 -1739 969
rect -1933 948 -1739 952
rect -1933 929 -1915 948
rect -1757 932 -1739 948
rect -841 968 -822 989
rect -747 968 -729 1568
rect -841 951 -729 968
rect -40 1570 -38 1576
rect -57 1540 -40 1559
rect -57 1504 -40 1523
rect -57 1434 -40 1487
rect -57 1346 -40 1417
rect -57 1269 -40 1329
rect -57 1187 -40 1252
rect -57 1107 -40 1170
rect -57 1050 -40 1090
rect -57 994 -40 1033
rect -841 930 -822 951
rect -57 944 -40 977
rect -57 893 -40 927
rect 928 894 958 905
rect -57 855 -40 876
rect 867 886 958 894
rect 867 869 877 886
rect 894 869 958 886
rect 867 861 958 869
rect 928 847 958 861
rect -2894 809 -2821 826
rect -1936 812 -1725 829
rect -840 812 -798 829
rect -57 813 -40 838
rect -99 779 -40 796
rect -3051 650 -3021 671
rect -2850 650 -2832 677
rect -1945 658 -1751 677
rect -3051 633 -2832 650
rect -3051 613 -3021 633
rect -2850 605 -2832 633
rect -2100 605 -2065 624
rect -99 607 -82 779
rect -51 739 -42 756
rect -25 739 12 756
rect -2211 452 -2157 460
rect -2211 435 -2193 452
rect -2176 435 -2157 452
rect -2211 421 -2157 435
rect -51 428 -17 441
rect -51 411 -42 428
rect -25 411 -17 428
rect -51 399 -17 411
rect -2105 310 -2073 329
rect -152 282 -17 327
rect -3052 174 -3022 189
rect -3052 145 -2817 174
rect -2083 160 -2051 169
rect -2083 157 -2076 160
rect -3052 131 -3022 145
rect -2187 143 -2076 157
rect -2059 143 -2051 160
rect -2187 122 -2051 143
rect -50 163 -17 282
rect -50 159 35 163
rect -50 134 114 159
rect -3052 31 -3022 52
rect -3052 14 -2849 31
rect -2101 14 -2066 33
rect 928 25 958 42
rect -3052 -6 -3022 14
rect 839 0 958 25
rect 928 -16 958 0
<< viali >>
rect -47 1595 -30 1612
rect -5 1595 12 1612
rect -1893 1322 -1874 1341
rect -1853 952 -1836 969
rect -57 1559 -40 1576
rect -57 1523 -40 1540
rect -57 1487 -40 1504
rect -57 1417 -40 1434
rect -57 1329 -40 1346
rect -57 1252 -40 1269
rect -57 1170 -40 1187
rect -57 1090 -40 1107
rect -57 1033 -40 1050
rect -57 977 -40 994
rect -57 927 -40 944
rect -57 876 -40 893
rect 877 869 894 886
rect -57 838 -40 855
rect -798 812 -781 829
rect -57 796 -40 813
rect -42 739 -25 756
rect -2193 435 -2176 452
rect -42 411 -25 428
rect -2076 143 -2059 160
<< metal1 >>
rect -61 1612 49 1616
rect -61 1595 -47 1612
rect -30 1595 -5 1612
rect 12 1595 49 1612
rect -61 1591 49 1595
rect -61 1576 -36 1591
rect -61 1559 -57 1576
rect -40 1559 -36 1576
rect -61 1540 -36 1559
rect -61 1523 -57 1540
rect -40 1523 -36 1540
rect -61 1504 -36 1523
rect -61 1487 -57 1504
rect -40 1487 -36 1504
rect -61 1434 -36 1487
rect -61 1417 -57 1434
rect -40 1417 -36 1434
rect -61 1346 -36 1417
rect -2678 1344 -1866 1345
rect -2923 1341 -1866 1344
rect -2923 1322 -1893 1341
rect -1874 1322 -1866 1341
rect -61 1329 -57 1346
rect -40 1329 -36 1346
rect -2923 1318 -1866 1322
rect -2923 229 -2897 1318
rect -1757 1278 -1723 1328
rect -61 1269 -36 1329
rect -61 1252 -57 1269
rect -40 1252 -36 1269
rect -61 1187 -36 1252
rect -61 1170 -57 1187
rect -40 1170 -36 1187
rect -61 1107 -36 1170
rect -61 1090 -57 1107
rect -40 1090 -36 1107
rect -61 1050 -36 1090
rect -61 1033 -57 1050
rect -40 1033 -36 1050
rect -1933 976 -1719 1008
rect -1933 947 -1859 976
rect -1829 947 -1719 976
rect -1933 912 -1719 947
rect -61 994 -36 1033
rect -61 977 -57 994
rect -40 977 -36 994
rect -61 944 -36 977
rect -61 927 -57 944
rect -40 927 -36 944
rect -61 893 -36 927
rect -61 876 -57 893
rect -40 876 -36 893
rect -61 855 -36 876
rect 860 891 909 894
rect 860 865 873 891
rect 899 865 909 891
rect 860 862 909 865
rect -61 838 -57 855
rect -40 838 -36 855
rect -806 834 -772 838
rect -806 808 -802 834
rect -776 808 -772 834
rect -806 804 -772 808
rect -61 813 -36 838
rect -61 802 -57 813
rect -103 796 -57 802
rect -40 796 -36 813
rect -103 777 -36 796
rect -2850 592 -2840 688
rect -2124 592 -2064 640
rect -103 624 -78 777
rect -51 756 -17 763
rect -51 730 -46 756
rect -20 730 -17 756
rect -51 727 -17 730
rect -2211 454 -2157 460
rect -2211 428 -2194 454
rect -2168 428 -2157 454
rect -2211 421 -2157 428
rect -51 433 -17 441
rect -51 407 -46 433
rect -20 407 -17 433
rect -51 402 -17 407
rect -2106 296 -2046 344
rect -2923 201 -2751 229
rect -2086 169 -2048 175
rect -2086 143 -2080 169
rect -2054 143 -2048 169
rect -2086 137 -2048 143
rect -2081 104 -2048 109
rect -2081 78 -2078 104
rect -2052 78 -2048 104
rect -2081 75 -2048 78
<< via1 >>
rect -1859 969 -1829 976
rect -1859 952 -1853 969
rect -1853 952 -1836 969
rect -1836 952 -1829 969
rect -1859 947 -1829 952
rect 873 886 899 891
rect 873 869 877 886
rect 877 869 894 886
rect 894 869 899 886
rect 873 865 899 869
rect -802 829 -776 834
rect -802 812 -798 829
rect -798 812 -781 829
rect -781 812 -776 829
rect -802 808 -776 812
rect -46 739 -42 756
rect -42 739 -25 756
rect -25 739 -20 756
rect -46 730 -20 739
rect -2194 452 -2168 454
rect -2194 435 -2193 452
rect -2193 435 -2176 452
rect -2176 435 -2168 452
rect -2194 428 -2168 435
rect -46 428 -20 433
rect -46 411 -42 428
rect -42 411 -25 428
rect -25 411 -20 428
rect -46 407 -20 411
rect -2080 160 -2054 169
rect -2080 143 -2076 160
rect -2076 143 -2059 160
rect -2059 143 -2054 160
rect -2078 78 -2052 104
<< metal2 >>
rect -3051 979 -3021 988
rect -2927 979 -1799 1008
rect -3051 976 -1799 979
rect -3051 947 -1859 976
rect -1829 947 -1799 976
rect -3051 939 -1799 947
rect -3051 930 -3021 939
rect -2927 912 -1799 939
rect -806 891 909 894
rect -806 865 873 891
rect 899 865 909 891
rect -806 861 909 865
rect -806 834 -772 861
rect -806 808 -802 834
rect -776 808 -772 834
rect -806 804 -772 808
rect -51 756 -17 763
rect -51 730 -46 756
rect -20 730 -17 756
rect -2197 454 -2165 457
rect -2197 428 -2194 454
rect -2168 428 -2165 454
rect -2197 344 -2165 428
rect -51 433 -17 730
rect -51 407 -46 433
rect -20 407 -17 433
rect -51 402 -17 407
rect -2256 308 -2165 344
rect -2256 114 -2220 308
rect -2083 169 -2048 272
rect -2083 143 -2080 169
rect -2054 143 -2048 169
rect -2083 137 -2048 143
rect -2256 104 -2041 114
rect -2256 78 -2078 104
rect -2052 78 -2041 104
rect -2256 68 -2041 78
use CP  CP_0
timestamp 1605998167
transform 1 0 -2083 0 1 0
box 0 0 2067 640
use VCO_new  VCO_new_0
timestamp 1633061951
transform 1 0 174 0 1 910
box -174 -910 721 844
use PFD  PFD_0
timestamp 1605977318
transform 1 0 -2850 0 1 0
box 0 0 767 640
use FD  FD_1
timestamp 1605926473
transform 1 0 -2850 0 1 960
box 0 0 935 320
use FD  FD_2
timestamp 1605926473
transform -1 0 -822 0 -1 960
box 0 0 935 320
use FD  FD_0
timestamp 1605926473
transform -1 0 -1915 0 -1 960
box 0 0 935 320
use FD  FD_3
timestamp 1605926473
transform 1 0 -1757 0 1 960
box 0 0 935 320
use FD  FD_4
timestamp 1605926473
transform -1 0 -822 0 -1 1600
box 0 0 935 320
<< labels >>
rlabel locali -3051 1404 -3051 1462 3 vdd#1
port 1 e
rlabel locali -3051 613 -3051 671 3 vdd#2
port 2 e
rlabel locali -3052 -6 -3052 52 3 vdd#3
port 3 e
rlabel metal2 -3051 930 -3051 988 3 gnd#1
port 4 e
rlabel locali 958 847 958 905 7 out
port 5 w
rlabel locali 958 -16 958 42 7 gnd#2
port 6 w
rlabel locali -3052 131 -3052 189 3 ref
port 7 e
<< end >>
