magic
tech sky130A
timestamp 1633061951
<< nwell >>
rect -47 653 662 826
rect -171 117 662 653
rect -47 -18 662 117
<< nmos >>
rect 0 -174 15 -66
rect 100 -174 115 -66
rect 200 -174 215 -66
rect 300 -174 315 -66
rect 400 -174 415 -66
rect 500 -174 515 -66
rect 600 -174 615 -66
rect -124 -701 -109 -201
rect -29 -245 471 -230
rect -29 -345 471 -330
rect 600 -333 615 -225
rect -29 -445 471 -430
rect -29 -545 471 -530
rect -29 -645 471 -630
rect -29 -745 471 -730
rect -29 -845 471 -830
<< pmos >>
rect -29 764 471 779
rect -29 664 471 679
rect -124 135 -109 635
rect -29 564 471 579
rect -29 464 471 479
rect -29 364 471 379
rect -29 264 471 279
rect -29 164 471 179
rect 600 159 615 579
rect 0 0 15 108
rect 100 0 115 108
rect 200 0 215 108
rect 300 0 315 108
rect 400 0 415 108
rect 500 0 515 108
rect 600 0 615 108
<< ndiff >>
rect -29 -74 0 -66
rect -29 -91 -23 -74
rect -6 -91 0 -74
rect -29 -111 0 -91
rect -29 -128 -23 -111
rect -6 -128 0 -111
rect -29 -149 0 -128
rect -29 -166 -23 -149
rect -6 -166 0 -149
rect -29 -174 0 -166
rect 15 -72 44 -66
rect 15 -89 21 -72
rect 38 -89 44 -72
rect 15 -111 44 -89
rect 15 -128 21 -111
rect 38 -128 44 -111
rect 15 -149 44 -128
rect 15 -166 21 -149
rect 38 -166 44 -149
rect 15 -174 44 -166
rect 71 -74 100 -66
rect 71 -91 77 -74
rect 94 -91 100 -74
rect 71 -111 100 -91
rect 71 -128 77 -111
rect 94 -128 100 -111
rect 71 -149 100 -128
rect 71 -166 77 -149
rect 94 -166 100 -149
rect 71 -174 100 -166
rect 115 -72 144 -66
rect 115 -89 121 -72
rect 138 -89 144 -72
rect 115 -112 144 -89
rect 115 -129 121 -112
rect 138 -129 144 -112
rect 115 -149 144 -129
rect 115 -166 121 -149
rect 138 -166 144 -149
rect 115 -174 144 -166
rect 171 -74 200 -66
rect 171 -91 177 -74
rect 194 -91 200 -74
rect 171 -111 200 -91
rect 171 -128 177 -111
rect 194 -128 200 -111
rect 171 -149 200 -128
rect 171 -166 177 -149
rect 194 -166 200 -149
rect 171 -174 200 -166
rect 215 -72 244 -66
rect 215 -89 221 -72
rect 238 -89 244 -72
rect 215 -112 244 -89
rect 215 -129 221 -112
rect 238 -129 244 -112
rect 215 -149 244 -129
rect 215 -166 221 -149
rect 238 -166 244 -149
rect 215 -174 244 -166
rect 271 -74 300 -66
rect 271 -91 277 -74
rect 294 -91 300 -74
rect 271 -111 300 -91
rect 271 -128 277 -111
rect 294 -128 300 -111
rect 271 -149 300 -128
rect 271 -166 277 -149
rect 294 -166 300 -149
rect 271 -174 300 -166
rect 315 -72 344 -66
rect 315 -89 321 -72
rect 338 -89 344 -72
rect 315 -111 344 -89
rect 315 -128 321 -111
rect 338 -128 344 -111
rect 315 -149 344 -128
rect 315 -166 321 -149
rect 338 -166 344 -149
rect 315 -174 344 -166
rect 371 -74 400 -66
rect 371 -91 377 -74
rect 394 -91 400 -74
rect 371 -111 400 -91
rect 371 -128 377 -111
rect 394 -128 400 -111
rect 371 -149 400 -128
rect 371 -166 377 -149
rect 394 -166 400 -149
rect 371 -174 400 -166
rect 415 -72 444 -66
rect 415 -89 421 -72
rect 438 -89 444 -72
rect 415 -111 444 -89
rect 415 -128 421 -111
rect 438 -128 444 -111
rect 415 -149 444 -128
rect 415 -166 421 -149
rect 438 -166 444 -149
rect 415 -174 444 -166
rect 471 -74 500 -66
rect 471 -91 477 -74
rect 494 -91 500 -74
rect 471 -111 500 -91
rect 471 -128 477 -111
rect 494 -128 500 -111
rect 471 -149 500 -128
rect 471 -166 477 -149
rect 494 -166 500 -149
rect 471 -174 500 -166
rect 515 -74 544 -66
rect 515 -91 521 -74
rect 538 -91 544 -74
rect 515 -111 544 -91
rect 515 -128 521 -111
rect 538 -128 544 -111
rect 515 -149 544 -128
rect 515 -166 521 -149
rect 538 -166 544 -149
rect 515 -174 544 -166
rect 571 -74 600 -66
rect 571 -91 577 -74
rect 594 -91 600 -74
rect 571 -111 600 -91
rect 571 -128 577 -111
rect 594 -128 600 -111
rect 571 -149 600 -128
rect 571 -166 577 -149
rect 594 -166 600 -149
rect 571 -174 600 -166
rect 615 -74 644 -66
rect 615 -91 621 -74
rect 638 -91 644 -74
rect 615 -111 644 -91
rect 615 -128 621 -111
rect 638 -128 644 -111
rect 615 -149 644 -128
rect 615 -166 621 -149
rect 638 -166 644 -149
rect 615 -174 644 -166
rect -153 -209 -124 -201
rect -153 -226 -147 -209
rect -130 -226 -124 -209
rect -153 -244 -124 -226
rect -153 -261 -147 -244
rect -130 -261 -124 -244
rect -153 -279 -124 -261
rect -153 -296 -147 -279
rect -130 -296 -124 -279
rect -153 -314 -124 -296
rect -153 -331 -147 -314
rect -130 -331 -124 -314
rect -153 -348 -124 -331
rect -153 -365 -147 -348
rect -130 -365 -124 -348
rect -153 -383 -124 -365
rect -153 -400 -147 -383
rect -130 -400 -124 -383
rect -153 -418 -124 -400
rect -153 -435 -147 -418
rect -130 -435 -124 -418
rect -153 -453 -124 -435
rect -153 -470 -147 -453
rect -130 -470 -124 -453
rect -153 -488 -124 -470
rect -153 -505 -147 -488
rect -130 -505 -124 -488
rect -153 -523 -124 -505
rect -153 -540 -147 -523
rect -130 -540 -124 -523
rect -153 -558 -124 -540
rect -153 -575 -147 -558
rect -130 -575 -124 -558
rect -153 -592 -124 -575
rect -153 -609 -147 -592
rect -130 -609 -124 -592
rect -153 -627 -124 -609
rect -153 -644 -147 -627
rect -130 -644 -124 -627
rect -153 -676 -124 -644
rect -153 -693 -147 -676
rect -130 -693 -124 -676
rect -153 -701 -124 -693
rect -109 -209 -80 -201
rect -109 -226 -103 -209
rect -86 -226 -80 -209
rect -109 -244 -80 -226
rect -109 -261 -103 -244
rect -86 -261 -80 -244
rect -109 -279 -80 -261
rect -109 -296 -103 -279
rect -86 -296 -80 -279
rect -109 -314 -80 -296
rect -109 -331 -103 -314
rect -86 -331 -80 -314
rect -109 -348 -80 -331
rect -109 -365 -103 -348
rect -86 -365 -80 -348
rect -109 -383 -80 -365
rect -109 -400 -103 -383
rect -86 -400 -80 -383
rect -109 -418 -80 -400
rect -109 -435 -103 -418
rect -86 -435 -80 -418
rect -109 -453 -80 -435
rect -109 -470 -103 -453
rect -86 -470 -80 -453
rect -109 -488 -80 -470
rect -109 -505 -103 -488
rect -86 -505 -80 -488
rect -109 -523 -80 -505
rect -109 -540 -103 -523
rect -86 -540 -80 -523
rect -109 -558 -80 -540
rect -109 -575 -103 -558
rect -86 -575 -80 -558
rect -109 -592 -80 -575
rect -109 -609 -103 -592
rect -86 -609 -80 -592
rect -109 -627 -80 -609
rect -109 -644 -103 -627
rect -86 -644 -80 -627
rect -109 -676 -80 -644
rect -109 -693 -103 -676
rect -86 -693 -80 -676
rect -109 -701 -80 -693
rect -29 -207 471 -201
rect -29 -224 -21 -207
rect -4 -224 56 -207
rect 73 -224 132 -207
rect 149 -224 209 -207
rect 226 -224 286 -207
rect 303 -224 362 -207
rect 379 -224 435 -207
rect 452 -224 471 -207
rect -29 -230 471 -224
rect 571 -233 600 -225
rect -29 -251 471 -245
rect -29 -268 -21 -251
rect -4 -268 24 -251
rect 41 -268 69 -251
rect 86 -268 113 -251
rect 130 -268 158 -251
rect 175 -268 203 -251
rect 220 -268 248 -251
rect 265 -268 293 -251
rect 310 -268 338 -251
rect 355 -268 383 -251
rect 400 -268 427 -251
rect 444 -268 471 -251
rect -29 -274 471 -268
rect 571 -250 577 -233
rect 594 -250 600 -233
rect 571 -271 600 -250
rect 571 -288 577 -271
rect 594 -288 600 -271
rect -29 -307 471 -301
rect -29 -324 -21 -307
rect -4 -324 24 -307
rect 41 -324 69 -307
rect 86 -324 114 -307
rect 131 -324 159 -307
rect 176 -324 204 -307
rect 221 -324 248 -307
rect 265 -324 293 -307
rect 310 -324 338 -307
rect 355 -324 383 -307
rect 400 -324 428 -307
rect 445 -324 471 -307
rect -29 -330 471 -324
rect 571 -308 600 -288
rect 571 -325 577 -308
rect 594 -325 600 -308
rect 571 -333 600 -325
rect 615 -233 644 -225
rect 615 -250 621 -233
rect 638 -250 644 -233
rect 615 -271 644 -250
rect 615 -288 621 -271
rect 638 -288 644 -271
rect 615 -308 644 -288
rect 615 -325 621 -308
rect 638 -325 644 -308
rect 615 -333 644 -325
rect -29 -351 471 -345
rect -29 -368 -21 -351
rect -4 -368 24 -351
rect 41 -368 69 -351
rect 86 -368 113 -351
rect 130 -368 158 -351
rect 175 -368 203 -351
rect 220 -368 248 -351
rect 265 -368 293 -351
rect 310 -368 338 -351
rect 355 -368 383 -351
rect 400 -368 427 -351
rect 444 -368 471 -351
rect -29 -374 471 -368
rect -29 -407 471 -401
rect -29 -424 -21 -407
rect -4 -424 24 -407
rect 41 -424 69 -407
rect 86 -424 114 -407
rect 131 -424 170 -407
rect 187 -424 209 -407
rect 226 -424 248 -407
rect 265 -424 288 -407
rect 305 -424 327 -407
rect 344 -424 366 -407
rect 383 -424 405 -407
rect 422 -424 444 -407
rect 461 -424 471 -407
rect -29 -430 471 -424
rect -29 -451 471 -445
rect -29 -468 -21 -451
rect -4 -468 18 -451
rect 35 -468 58 -451
rect 75 -468 97 -451
rect 114 -468 136 -451
rect 153 -468 175 -451
rect 192 -468 214 -451
rect 231 -468 254 -451
rect 271 -468 293 -451
rect 310 -468 332 -451
rect 349 -468 371 -451
rect 388 -468 411 -451
rect 428 -468 445 -451
rect 462 -468 471 -451
rect -29 -474 471 -468
rect -29 -507 471 -501
rect -29 -524 -21 -507
rect -4 -524 18 -507
rect 35 -524 58 -507
rect 75 -524 97 -507
rect 114 -524 136 -507
rect 153 -524 175 -507
rect 192 -524 214 -507
rect 231 -524 254 -507
rect 271 -524 288 -507
rect 305 -524 327 -507
rect 344 -524 366 -507
rect 383 -524 406 -507
rect 423 -524 445 -507
rect 462 -524 471 -507
rect -29 -530 471 -524
rect -29 -551 471 -545
rect -29 -568 -21 -551
rect -4 -568 24 -551
rect 41 -568 69 -551
rect 86 -568 113 -551
rect 130 -568 158 -551
rect 175 -568 203 -551
rect 220 -568 248 -551
rect 265 -568 293 -551
rect 310 -568 338 -551
rect 355 -568 383 -551
rect 400 -568 427 -551
rect 444 -568 471 -551
rect -29 -574 471 -568
rect -29 -607 471 -601
rect -29 -624 -21 -607
rect -4 -624 24 -607
rect 41 -624 69 -607
rect 86 -624 114 -607
rect 131 -624 158 -607
rect 175 -624 203 -607
rect 220 -624 248 -607
rect 265 -624 293 -607
rect 310 -624 338 -607
rect 355 -624 383 -607
rect 400 -624 428 -607
rect 445 -624 471 -607
rect -29 -630 471 -624
rect -29 -651 471 -645
rect -29 -668 -21 -651
rect -4 -668 29 -651
rect 46 -668 80 -651
rect 97 -668 130 -651
rect 147 -668 181 -651
rect 198 -668 231 -651
rect 248 -668 282 -651
rect 299 -668 332 -651
rect 349 -668 383 -651
rect 400 -668 428 -651
rect 445 -668 471 -651
rect -29 -674 471 -668
rect -29 -707 471 -701
rect -29 -724 -21 -707
rect -4 -724 24 -707
rect 41 -724 69 -707
rect 86 -724 114 -707
rect 131 -724 158 -707
rect 175 -724 203 -707
rect 220 -724 248 -707
rect 265 -724 293 -707
rect 310 -724 338 -707
rect 355 -724 383 -707
rect 400 -724 428 -707
rect 445 -724 471 -707
rect -29 -730 471 -724
rect -29 -751 471 -745
rect -29 -768 -21 -751
rect -4 -768 24 -751
rect 41 -768 69 -751
rect 86 -768 113 -751
rect 130 -768 158 -751
rect 175 -768 203 -751
rect 220 -768 248 -751
rect 265 -768 293 -751
rect 310 -768 338 -751
rect 355 -768 373 -751
rect 390 -768 427 -751
rect 444 -768 471 -751
rect -29 -774 471 -768
rect -29 -807 471 -801
rect -29 -824 -21 -807
rect -4 -824 24 -807
rect 41 -824 69 -807
rect 86 -824 113 -807
rect 130 -824 158 -807
rect 175 -824 203 -807
rect 220 -824 248 -807
rect 265 -824 293 -807
rect 310 -824 338 -807
rect 355 -824 383 -807
rect 400 -824 427 -807
rect 444 -824 471 -807
rect -29 -830 471 -824
rect -29 -851 471 -845
rect -29 -868 -21 -851
rect -4 -868 24 -851
rect 41 -868 63 -851
rect 80 -868 102 -851
rect 119 -868 147 -851
rect 164 -868 192 -851
rect 209 -868 237 -851
rect 254 -868 282 -851
rect 299 -868 327 -851
rect 344 -868 371 -851
rect 388 -868 416 -851
rect 433 -868 450 -851
rect 467 -868 471 -851
rect -29 -874 471 -868
<< pdiff >>
rect -29 802 471 808
rect -29 785 -21 802
rect -4 785 38 802
rect 55 785 98 802
rect 115 785 157 802
rect 174 785 216 802
rect 233 785 276 802
rect 293 785 335 802
rect 352 785 394 802
rect 411 785 439 802
rect 456 785 471 802
rect -29 779 471 785
rect -29 758 471 764
rect -29 741 -21 758
rect -4 741 46 758
rect 63 741 113 758
rect 130 741 180 758
rect 197 741 247 758
rect 264 741 315 758
rect 332 741 382 758
rect 399 741 425 758
rect 442 741 471 758
rect -29 735 471 741
rect -29 702 471 708
rect -29 685 -21 702
rect -4 685 38 702
rect 55 685 98 702
rect 115 685 157 702
rect 174 685 216 702
rect 233 685 276 702
rect 293 685 335 702
rect 352 685 394 702
rect 411 685 439 702
rect 456 685 471 702
rect -29 679 471 685
rect -153 627 -124 635
rect -153 610 -147 627
rect -130 610 -124 627
rect -153 592 -124 610
rect -153 575 -147 592
rect -130 575 -124 592
rect -153 549 -124 575
rect -153 532 -147 549
rect -130 532 -124 549
rect -153 507 -124 532
rect -153 490 -147 507
rect -130 490 -124 507
rect -153 464 -124 490
rect -153 447 -147 464
rect -130 447 -124 464
rect -153 422 -124 447
rect -153 405 -147 422
rect -130 405 -124 422
rect -153 379 -124 405
rect -153 362 -147 379
rect -130 362 -124 379
rect -153 337 -124 362
rect -153 320 -147 337
rect -130 320 -124 337
rect -153 294 -124 320
rect -153 277 -147 294
rect -130 277 -124 294
rect -153 252 -124 277
rect -153 235 -147 252
rect -130 235 -124 252
rect -153 209 -124 235
rect -153 192 -147 209
rect -130 192 -124 209
rect -153 160 -124 192
rect -153 143 -147 160
rect -130 143 -124 160
rect -153 135 -124 143
rect -109 627 -80 635
rect -109 610 -103 627
rect -86 610 -80 627
rect -109 592 -80 610
rect -109 575 -103 592
rect -86 575 -80 592
rect -109 549 -80 575
rect -109 532 -103 549
rect -86 532 -80 549
rect -109 507 -80 532
rect -109 490 -103 507
rect -86 490 -80 507
rect -109 464 -80 490
rect -109 447 -103 464
rect -86 447 -80 464
rect -109 422 -80 447
rect -109 405 -103 422
rect -86 405 -80 422
rect -109 379 -80 405
rect -109 362 -103 379
rect -86 362 -80 379
rect -109 337 -80 362
rect -109 320 -103 337
rect -86 320 -80 337
rect -109 294 -80 320
rect -109 277 -103 294
rect -86 277 -80 294
rect -109 252 -80 277
rect -109 235 -103 252
rect -86 235 -80 252
rect -109 209 -80 235
rect -109 192 -103 209
rect -86 192 -80 209
rect -109 160 -80 192
rect -109 143 -103 160
rect -86 143 -80 160
rect -109 135 -80 143
rect -29 658 471 664
rect -29 641 -21 658
rect -4 641 26 658
rect 43 641 64 658
rect 81 641 111 658
rect 128 641 158 658
rect 175 641 195 658
rect 212 641 243 658
rect 260 641 287 658
rect 304 641 327 658
rect 344 641 374 658
rect 391 641 433 658
rect 450 641 471 658
rect -29 635 471 641
rect -29 602 471 608
rect -29 585 -21 602
rect -4 585 38 602
rect 55 585 98 602
rect 115 585 157 602
rect 174 585 216 602
rect 233 585 276 602
rect 293 585 335 602
rect 352 585 394 602
rect 411 585 439 602
rect 456 585 471 602
rect -29 579 471 585
rect 571 571 600 579
rect -29 558 471 564
rect -29 541 -21 558
rect -4 541 19 558
rect 36 541 75 558
rect 92 541 122 558
rect 139 541 171 558
rect 188 541 224 558
rect 241 541 268 558
rect 285 541 312 558
rect 329 541 364 558
rect 381 541 445 558
rect 462 541 471 558
rect -29 535 471 541
rect 571 554 577 571
rect 594 554 600 571
rect 571 531 600 554
rect 571 514 577 531
rect 594 514 600 531
rect -29 502 471 508
rect -29 485 -21 502
rect -4 485 38 502
rect 55 485 98 502
rect 115 485 157 502
rect 174 485 216 502
rect 233 485 276 502
rect 293 485 335 502
rect 352 485 394 502
rect 411 485 439 502
rect 456 485 471 502
rect -29 479 471 485
rect 571 491 600 514
rect 571 474 577 491
rect 594 474 600 491
rect -29 458 471 464
rect -29 441 -21 458
rect -4 441 32 458
rect 49 441 89 458
rect 106 441 134 458
rect 151 441 199 458
rect 216 441 237 458
rect 254 441 285 458
rect 302 441 329 458
rect 346 441 381 458
rect 398 441 442 458
rect 459 441 471 458
rect -29 435 471 441
rect 571 452 600 474
rect 571 435 577 452
rect 594 435 600 452
rect 571 412 600 435
rect -29 402 471 408
rect -29 385 -21 402
rect -4 385 38 402
rect 55 385 98 402
rect 115 385 157 402
rect 174 385 216 402
rect 233 385 276 402
rect 293 385 335 402
rect 352 385 394 402
rect 411 385 439 402
rect 456 385 471 402
rect -29 379 471 385
rect 571 395 577 412
rect 594 395 600 412
rect 571 372 600 395
rect -29 358 471 364
rect -29 341 -21 358
rect -4 341 16 358
rect 33 341 75 358
rect 92 341 119 358
rect 136 341 171 358
rect 188 341 221 358
rect 238 341 267 358
rect 284 341 324 358
rect 341 341 363 358
rect 380 341 412 358
rect 429 341 446 358
rect 463 341 471 358
rect -29 335 471 341
rect 571 355 577 372
rect 594 355 600 372
rect 571 332 600 355
rect 571 315 577 332
rect 594 315 600 332
rect -29 302 471 308
rect -29 285 -21 302
rect -4 285 38 302
rect 55 285 98 302
rect 115 285 157 302
rect 174 285 216 302
rect 233 285 276 302
rect 293 285 335 302
rect 352 285 394 302
rect 411 285 439 302
rect 456 285 471 302
rect -29 279 471 285
rect 571 293 600 315
rect 571 276 577 293
rect 594 276 600 293
rect -29 258 471 264
rect -29 241 -21 258
rect -4 241 27 258
rect 44 241 86 258
rect 103 241 160 258
rect 177 241 234 258
rect 251 241 299 258
rect 316 241 363 258
rect 380 241 428 258
rect 445 241 471 258
rect -29 235 471 241
rect 571 253 600 276
rect 571 236 577 253
rect 594 236 600 253
rect 571 218 600 236
rect -29 202 471 208
rect -29 185 -21 202
rect -4 185 38 202
rect 55 185 98 202
rect 115 185 157 202
rect 174 185 216 202
rect 233 185 276 202
rect 293 185 335 202
rect 352 185 394 202
rect 411 185 439 202
rect 456 185 471 202
rect -29 179 471 185
rect 571 201 577 218
rect 594 201 600 218
rect 571 184 600 201
rect 571 167 577 184
rect 594 167 600 184
rect -29 158 471 164
rect 571 159 600 167
rect 615 571 644 579
rect 615 554 621 571
rect 638 554 644 571
rect 615 531 644 554
rect 615 514 621 531
rect 638 514 644 531
rect 615 491 644 514
rect 615 474 621 491
rect 638 474 644 491
rect 615 452 644 474
rect 615 435 621 452
rect 638 435 644 452
rect 615 412 644 435
rect 615 395 621 412
rect 638 395 644 412
rect 615 372 644 395
rect 615 355 621 372
rect 638 355 644 372
rect 615 332 644 355
rect 615 315 621 332
rect 638 315 644 332
rect 615 293 644 315
rect 615 276 621 293
rect 638 276 644 293
rect 615 253 644 276
rect 615 236 621 253
rect 638 236 644 253
rect 615 218 644 236
rect 615 201 621 218
rect 638 201 644 218
rect 615 184 644 201
rect 615 167 621 184
rect 638 167 644 184
rect 615 159 644 167
rect -29 141 -21 158
rect -4 141 36 158
rect 53 141 93 158
rect 110 141 150 158
rect 167 141 207 158
rect 224 141 264 158
rect 281 141 321 158
rect 338 141 378 158
rect 395 141 435 158
rect 452 141 471 158
rect -29 135 471 141
rect -29 100 0 108
rect -29 83 -23 100
rect -6 83 0 100
rect -29 63 0 83
rect -29 46 -23 63
rect -6 46 0 63
rect -29 25 0 46
rect -29 8 -23 25
rect -6 8 0 25
rect -29 0 0 8
rect 15 100 44 108
rect 15 83 21 100
rect 38 83 44 100
rect 15 63 44 83
rect 15 46 21 63
rect 38 46 44 63
rect 15 23 44 46
rect 15 6 21 23
rect 38 6 44 23
rect 15 0 44 6
rect 71 100 100 108
rect 71 83 77 100
rect 94 83 100 100
rect 71 66 100 83
rect 71 49 77 66
rect 94 49 100 66
rect 71 25 100 49
rect 71 8 77 25
rect 94 8 100 25
rect 71 0 100 8
rect 115 100 144 108
rect 115 83 121 100
rect 138 83 144 100
rect 115 63 144 83
rect 115 46 121 63
rect 138 46 144 63
rect 115 23 144 46
rect 115 6 121 23
rect 138 6 144 23
rect 115 0 144 6
rect 171 100 200 108
rect 171 83 177 100
rect 194 83 200 100
rect 171 66 200 83
rect 171 49 177 66
rect 194 49 200 66
rect 171 25 200 49
rect 171 8 177 25
rect 194 8 200 25
rect 171 0 200 8
rect 215 100 244 108
rect 215 83 221 100
rect 238 83 244 100
rect 215 63 244 83
rect 215 46 221 63
rect 238 46 244 63
rect 215 23 244 46
rect 215 6 221 23
rect 238 6 244 23
rect 215 0 244 6
rect 271 100 300 108
rect 271 83 277 100
rect 294 83 300 100
rect 271 66 300 83
rect 271 49 277 66
rect 294 49 300 66
rect 271 25 300 49
rect 271 8 277 25
rect 294 8 300 25
rect 271 0 300 8
rect 315 100 344 108
rect 315 83 321 100
rect 338 83 344 100
rect 315 63 344 83
rect 315 46 321 63
rect 338 46 344 63
rect 315 23 344 46
rect 315 6 321 23
rect 338 6 344 23
rect 315 0 344 6
rect 371 100 400 108
rect 371 83 377 100
rect 394 83 400 100
rect 371 66 400 83
rect 371 49 377 66
rect 394 49 400 66
rect 371 25 400 49
rect 371 8 377 25
rect 394 8 400 25
rect 371 0 400 8
rect 415 100 444 108
rect 415 83 421 100
rect 438 83 444 100
rect 415 63 444 83
rect 415 46 421 63
rect 438 46 444 63
rect 415 23 444 46
rect 415 6 421 23
rect 438 6 444 23
rect 415 0 444 6
rect 471 100 500 108
rect 471 83 477 100
rect 494 83 500 100
rect 471 66 500 83
rect 471 49 477 66
rect 494 49 500 66
rect 471 25 500 49
rect 471 8 477 25
rect 494 8 500 25
rect 471 0 500 8
rect 515 100 544 108
rect 515 83 521 100
rect 538 83 544 100
rect 515 66 544 83
rect 515 49 521 66
rect 538 49 544 66
rect 515 23 544 49
rect 515 6 521 23
rect 538 6 544 23
rect 515 0 544 6
rect 571 100 600 108
rect 571 83 577 100
rect 594 83 600 100
rect 571 66 600 83
rect 571 49 577 66
rect 594 49 600 66
rect 571 25 600 49
rect 571 8 577 25
rect 594 8 600 25
rect 571 0 600 8
rect 615 100 644 108
rect 615 83 621 100
rect 638 83 644 100
rect 615 66 644 83
rect 615 49 621 66
rect 638 49 644 66
rect 615 23 644 49
rect 615 6 621 23
rect 638 6 644 23
rect 615 0 644 6
<< ndiffc >>
rect -23 -91 -6 -74
rect -23 -128 -6 -111
rect -23 -166 -6 -149
rect 21 -89 38 -72
rect 21 -128 38 -111
rect 21 -166 38 -149
rect 77 -91 94 -74
rect 77 -128 94 -111
rect 77 -166 94 -149
rect 121 -89 138 -72
rect 121 -129 138 -112
rect 121 -166 138 -149
rect 177 -91 194 -74
rect 177 -128 194 -111
rect 177 -166 194 -149
rect 221 -89 238 -72
rect 221 -129 238 -112
rect 221 -166 238 -149
rect 277 -91 294 -74
rect 277 -128 294 -111
rect 277 -166 294 -149
rect 321 -89 338 -72
rect 321 -128 338 -111
rect 321 -166 338 -149
rect 377 -91 394 -74
rect 377 -128 394 -111
rect 377 -166 394 -149
rect 421 -89 438 -72
rect 421 -128 438 -111
rect 421 -166 438 -149
rect 477 -91 494 -74
rect 477 -128 494 -111
rect 477 -166 494 -149
rect 521 -91 538 -74
rect 521 -128 538 -111
rect 521 -166 538 -149
rect 577 -91 594 -74
rect 577 -128 594 -111
rect 577 -166 594 -149
rect 621 -91 638 -74
rect 621 -128 638 -111
rect 621 -166 638 -149
rect -147 -226 -130 -209
rect -147 -261 -130 -244
rect -147 -296 -130 -279
rect -147 -331 -130 -314
rect -147 -365 -130 -348
rect -147 -400 -130 -383
rect -147 -435 -130 -418
rect -147 -470 -130 -453
rect -147 -505 -130 -488
rect -147 -540 -130 -523
rect -147 -575 -130 -558
rect -147 -609 -130 -592
rect -147 -644 -130 -627
rect -147 -693 -130 -676
rect -103 -226 -86 -209
rect -103 -261 -86 -244
rect -103 -296 -86 -279
rect -103 -331 -86 -314
rect -103 -365 -86 -348
rect -103 -400 -86 -383
rect -103 -435 -86 -418
rect -103 -470 -86 -453
rect -103 -505 -86 -488
rect -103 -540 -86 -523
rect -103 -575 -86 -558
rect -103 -609 -86 -592
rect -103 -644 -86 -627
rect -103 -693 -86 -676
rect -21 -224 -4 -207
rect 56 -224 73 -207
rect 132 -224 149 -207
rect 209 -224 226 -207
rect 286 -224 303 -207
rect 362 -224 379 -207
rect 435 -224 452 -207
rect -21 -268 -4 -251
rect 24 -268 41 -251
rect 69 -268 86 -251
rect 113 -268 130 -251
rect 158 -268 175 -251
rect 203 -268 220 -251
rect 248 -268 265 -251
rect 293 -268 310 -251
rect 338 -268 355 -251
rect 383 -268 400 -251
rect 427 -268 444 -251
rect 577 -250 594 -233
rect 577 -288 594 -271
rect -21 -324 -4 -307
rect 24 -324 41 -307
rect 69 -324 86 -307
rect 114 -324 131 -307
rect 159 -324 176 -307
rect 204 -324 221 -307
rect 248 -324 265 -307
rect 293 -324 310 -307
rect 338 -324 355 -307
rect 383 -324 400 -307
rect 428 -324 445 -307
rect 577 -325 594 -308
rect 621 -250 638 -233
rect 621 -288 638 -271
rect 621 -325 638 -308
rect -21 -368 -4 -351
rect 24 -368 41 -351
rect 69 -368 86 -351
rect 113 -368 130 -351
rect 158 -368 175 -351
rect 203 -368 220 -351
rect 248 -368 265 -351
rect 293 -368 310 -351
rect 338 -368 355 -351
rect 383 -368 400 -351
rect 427 -368 444 -351
rect -21 -424 -4 -407
rect 24 -424 41 -407
rect 69 -424 86 -407
rect 114 -424 131 -407
rect 170 -424 187 -407
rect 209 -424 226 -407
rect 248 -424 265 -407
rect 288 -424 305 -407
rect 327 -424 344 -407
rect 366 -424 383 -407
rect 405 -424 422 -407
rect 444 -424 461 -407
rect -21 -468 -4 -451
rect 18 -468 35 -451
rect 58 -468 75 -451
rect 97 -468 114 -451
rect 136 -468 153 -451
rect 175 -468 192 -451
rect 214 -468 231 -451
rect 254 -468 271 -451
rect 293 -468 310 -451
rect 332 -468 349 -451
rect 371 -468 388 -451
rect 411 -468 428 -451
rect 445 -468 462 -451
rect -21 -524 -4 -507
rect 18 -524 35 -507
rect 58 -524 75 -507
rect 97 -524 114 -507
rect 136 -524 153 -507
rect 175 -524 192 -507
rect 214 -524 231 -507
rect 254 -524 271 -507
rect 288 -524 305 -507
rect 327 -524 344 -507
rect 366 -524 383 -507
rect 406 -524 423 -507
rect 445 -524 462 -507
rect -21 -568 -4 -551
rect 24 -568 41 -551
rect 69 -568 86 -551
rect 113 -568 130 -551
rect 158 -568 175 -551
rect 203 -568 220 -551
rect 248 -568 265 -551
rect 293 -568 310 -551
rect 338 -568 355 -551
rect 383 -568 400 -551
rect 427 -568 444 -551
rect -21 -624 -4 -607
rect 24 -624 41 -607
rect 69 -624 86 -607
rect 114 -624 131 -607
rect 158 -624 175 -607
rect 203 -624 220 -607
rect 248 -624 265 -607
rect 293 -624 310 -607
rect 338 -624 355 -607
rect 383 -624 400 -607
rect 428 -624 445 -607
rect -21 -668 -4 -651
rect 29 -668 46 -651
rect 80 -668 97 -651
rect 130 -668 147 -651
rect 181 -668 198 -651
rect 231 -668 248 -651
rect 282 -668 299 -651
rect 332 -668 349 -651
rect 383 -668 400 -651
rect 428 -668 445 -651
rect -21 -724 -4 -707
rect 24 -724 41 -707
rect 69 -724 86 -707
rect 114 -724 131 -707
rect 158 -724 175 -707
rect 203 -724 220 -707
rect 248 -724 265 -707
rect 293 -724 310 -707
rect 338 -724 355 -707
rect 383 -724 400 -707
rect 428 -724 445 -707
rect -21 -768 -4 -751
rect 24 -768 41 -751
rect 69 -768 86 -751
rect 113 -768 130 -751
rect 158 -768 175 -751
rect 203 -768 220 -751
rect 248 -768 265 -751
rect 293 -768 310 -751
rect 338 -768 355 -751
rect 373 -768 390 -751
rect 427 -768 444 -751
rect -21 -824 -4 -807
rect 24 -824 41 -807
rect 69 -824 86 -807
rect 113 -824 130 -807
rect 158 -824 175 -807
rect 203 -824 220 -807
rect 248 -824 265 -807
rect 293 -824 310 -807
rect 338 -824 355 -807
rect 383 -824 400 -807
rect 427 -824 444 -807
rect -21 -868 -4 -851
rect 24 -868 41 -851
rect 63 -868 80 -851
rect 102 -868 119 -851
rect 147 -868 164 -851
rect 192 -868 209 -851
rect 237 -868 254 -851
rect 282 -868 299 -851
rect 327 -868 344 -851
rect 371 -868 388 -851
rect 416 -868 433 -851
rect 450 -868 467 -851
<< pdiffc >>
rect -21 785 -4 802
rect 38 785 55 802
rect 98 785 115 802
rect 157 785 174 802
rect 216 785 233 802
rect 276 785 293 802
rect 335 785 352 802
rect 394 785 411 802
rect 439 785 456 802
rect -21 741 -4 758
rect 46 741 63 758
rect 113 741 130 758
rect 180 741 197 758
rect 247 741 264 758
rect 315 741 332 758
rect 382 741 399 758
rect 425 741 442 758
rect -21 685 -4 702
rect 38 685 55 702
rect 98 685 115 702
rect 157 685 174 702
rect 216 685 233 702
rect 276 685 293 702
rect 335 685 352 702
rect 394 685 411 702
rect 439 685 456 702
rect -147 610 -130 627
rect -147 575 -130 592
rect -147 532 -130 549
rect -147 490 -130 507
rect -147 447 -130 464
rect -147 405 -130 422
rect -147 362 -130 379
rect -147 320 -130 337
rect -147 277 -130 294
rect -147 235 -130 252
rect -147 192 -130 209
rect -147 143 -130 160
rect -103 610 -86 627
rect -103 575 -86 592
rect -103 532 -86 549
rect -103 490 -86 507
rect -103 447 -86 464
rect -103 405 -86 422
rect -103 362 -86 379
rect -103 320 -86 337
rect -103 277 -86 294
rect -103 235 -86 252
rect -103 192 -86 209
rect -103 143 -86 160
rect -21 641 -4 658
rect 26 641 43 658
rect 64 641 81 658
rect 111 641 128 658
rect 158 641 175 658
rect 195 641 212 658
rect 243 641 260 658
rect 287 641 304 658
rect 327 641 344 658
rect 374 641 391 658
rect 433 641 450 658
rect -21 585 -4 602
rect 38 585 55 602
rect 98 585 115 602
rect 157 585 174 602
rect 216 585 233 602
rect 276 585 293 602
rect 335 585 352 602
rect 394 585 411 602
rect 439 585 456 602
rect -21 541 -4 558
rect 19 541 36 558
rect 75 541 92 558
rect 122 541 139 558
rect 171 541 188 558
rect 224 541 241 558
rect 268 541 285 558
rect 312 541 329 558
rect 364 541 381 558
rect 445 541 462 558
rect 577 554 594 571
rect 577 514 594 531
rect -21 485 -4 502
rect 38 485 55 502
rect 98 485 115 502
rect 157 485 174 502
rect 216 485 233 502
rect 276 485 293 502
rect 335 485 352 502
rect 394 485 411 502
rect 439 485 456 502
rect 577 474 594 491
rect -21 441 -4 458
rect 32 441 49 458
rect 89 441 106 458
rect 134 441 151 458
rect 199 441 216 458
rect 237 441 254 458
rect 285 441 302 458
rect 329 441 346 458
rect 381 441 398 458
rect 442 441 459 458
rect 577 435 594 452
rect -21 385 -4 402
rect 38 385 55 402
rect 98 385 115 402
rect 157 385 174 402
rect 216 385 233 402
rect 276 385 293 402
rect 335 385 352 402
rect 394 385 411 402
rect 439 385 456 402
rect 577 395 594 412
rect -21 341 -4 358
rect 16 341 33 358
rect 75 341 92 358
rect 119 341 136 358
rect 171 341 188 358
rect 221 341 238 358
rect 267 341 284 358
rect 324 341 341 358
rect 363 341 380 358
rect 412 341 429 358
rect 446 341 463 358
rect 577 355 594 372
rect 577 315 594 332
rect -21 285 -4 302
rect 38 285 55 302
rect 98 285 115 302
rect 157 285 174 302
rect 216 285 233 302
rect 276 285 293 302
rect 335 285 352 302
rect 394 285 411 302
rect 439 285 456 302
rect 577 276 594 293
rect -21 241 -4 258
rect 27 241 44 258
rect 86 241 103 258
rect 160 241 177 258
rect 234 241 251 258
rect 299 241 316 258
rect 363 241 380 258
rect 428 241 445 258
rect 577 236 594 253
rect -21 185 -4 202
rect 38 185 55 202
rect 98 185 115 202
rect 157 185 174 202
rect 216 185 233 202
rect 276 185 293 202
rect 335 185 352 202
rect 394 185 411 202
rect 439 185 456 202
rect 577 201 594 218
rect 577 167 594 184
rect 621 554 638 571
rect 621 514 638 531
rect 621 474 638 491
rect 621 435 638 452
rect 621 395 638 412
rect 621 355 638 372
rect 621 315 638 332
rect 621 276 638 293
rect 621 236 638 253
rect 621 201 638 218
rect 621 167 638 184
rect -21 141 -4 158
rect 36 141 53 158
rect 93 141 110 158
rect 150 141 167 158
rect 207 141 224 158
rect 264 141 281 158
rect 321 141 338 158
rect 378 141 395 158
rect 435 141 452 158
rect -23 83 -6 100
rect -23 46 -6 63
rect -23 8 -6 25
rect 21 83 38 100
rect 21 46 38 63
rect 21 6 38 23
rect 77 83 94 100
rect 77 49 94 66
rect 77 8 94 25
rect 121 83 138 100
rect 121 46 138 63
rect 121 6 138 23
rect 177 83 194 100
rect 177 49 194 66
rect 177 8 194 25
rect 221 83 238 100
rect 221 46 238 63
rect 221 6 238 23
rect 277 83 294 100
rect 277 49 294 66
rect 277 8 294 25
rect 321 83 338 100
rect 321 46 338 63
rect 321 6 338 23
rect 377 83 394 100
rect 377 49 394 66
rect 377 8 394 25
rect 421 83 438 100
rect 421 46 438 63
rect 421 6 438 23
rect 477 83 494 100
rect 477 49 494 66
rect 477 8 494 25
rect 521 83 538 100
rect 521 49 538 66
rect 521 6 538 23
rect 577 83 594 100
rect 577 49 594 66
rect 577 8 594 25
rect 621 83 638 100
rect 621 49 638 66
rect 621 6 638 23
<< poly >>
rect -52 764 -29 779
rect 471 764 484 779
rect -52 679 -37 764
rect -52 664 -29 679
rect 471 664 484 679
rect -124 635 -109 648
rect -52 579 -37 664
rect 600 587 669 602
rect 600 579 615 587
rect -52 564 -29 579
rect 471 564 484 579
rect -52 479 -37 564
rect -52 464 -29 479
rect 471 464 484 479
rect -52 379 -37 464
rect -52 364 -29 379
rect 471 364 484 379
rect -52 279 -37 364
rect -52 264 -29 279
rect 471 264 484 279
rect -52 179 -37 264
rect -52 164 -29 179
rect 471 164 484 179
rect -124 117 -109 135
rect -52 117 -37 164
rect 600 146 615 159
rect -124 110 -37 117
rect -124 93 -103 110
rect -86 93 -37 110
rect 0 108 15 121
rect 100 108 115 121
rect 200 108 215 121
rect 300 108 315 121
rect 400 108 415 121
rect 500 108 515 121
rect 600 108 615 121
rect -124 86 -37 93
rect 0 -18 15 0
rect 100 -18 115 0
rect 200 -18 215 0
rect 300 -18 315 0
rect 400 -18 415 0
rect 500 -18 515 0
rect 600 -18 615 0
rect 652 -16 669 587
rect -29 -25 15 -18
rect -29 -42 -21 -25
rect -4 -42 15 -25
rect -29 -49 15 -42
rect 71 -25 115 -18
rect 71 -42 79 -25
rect 96 -42 115 -25
rect 71 -49 115 -42
rect 171 -25 215 -18
rect 171 -42 179 -25
rect 196 -42 215 -25
rect 171 -49 215 -42
rect 271 -25 315 -18
rect 271 -42 279 -25
rect 296 -42 315 -25
rect 271 -49 315 -42
rect 371 -25 415 -18
rect 371 -42 379 -25
rect 396 -42 415 -25
rect 371 -49 415 -42
rect 471 -25 515 -18
rect 471 -42 479 -25
rect 496 -42 515 -25
rect 471 -49 515 -42
rect 571 -25 615 -18
rect 571 -42 579 -25
rect 596 -42 615 -25
rect 571 -49 615 -42
rect 636 -24 669 -16
rect 636 -41 644 -24
rect 661 -41 669 -24
rect 636 -49 669 -41
rect 0 -66 15 -49
rect 100 -66 115 -49
rect 200 -66 215 -49
rect 300 -66 315 -49
rect 400 -66 415 -49
rect 500 -66 515 -49
rect 600 -66 615 -49
rect -166 -154 -37 -147
rect -166 -171 -158 -154
rect -141 -171 -37 -154
rect -166 -178 -37 -171
rect -124 -201 -109 -178
rect -52 -230 -37 -178
rect 0 -187 15 -174
rect 100 -187 115 -174
rect 200 -187 215 -174
rect 300 -187 315 -174
rect 400 -187 415 -174
rect 500 -187 515 -174
rect 600 -187 615 -174
rect 600 -225 615 -212
rect -52 -245 -29 -230
rect 471 -245 484 -230
rect -52 -330 -37 -245
rect -52 -345 -29 -330
rect 471 -345 484 -330
rect 600 -341 615 -333
rect 652 -341 669 -49
rect -52 -430 -37 -345
rect 600 -356 669 -341
rect -52 -445 -29 -430
rect 471 -445 484 -430
rect -52 -530 -37 -445
rect -52 -545 -29 -530
rect 471 -545 484 -530
rect -52 -630 -37 -545
rect -52 -645 -29 -630
rect 471 -645 484 -630
rect -124 -714 -109 -701
rect -52 -730 -37 -645
rect -52 -745 -29 -730
rect 471 -745 484 -730
rect -52 -830 -37 -745
rect -52 -845 -29 -830
rect 471 -845 484 -830
<< polycont >>
rect -103 93 -86 110
rect -21 -42 -4 -25
rect 79 -42 96 -25
rect 179 -42 196 -25
rect 279 -42 296 -25
rect 379 -42 396 -25
rect 479 -42 496 -25
rect 579 -42 596 -25
rect 644 -41 661 -24
rect -158 -171 -141 -154
<< locali >>
rect -63 840 670 844
rect -63 823 -55 840
rect -38 823 -18 840
rect -1 823 26 840
rect 43 823 71 840
rect 88 823 115 840
rect 132 823 159 840
rect 176 823 204 840
rect 221 823 248 840
rect 265 823 292 840
rect 309 823 336 840
rect 353 823 381 840
rect 398 823 425 840
rect 442 823 469 840
rect 486 823 514 840
rect 531 823 558 840
rect 575 823 602 840
rect 619 823 647 840
rect 664 823 670 840
rect -63 819 670 823
rect -63 798 -46 819
rect -29 785 -21 802
rect -4 785 38 802
rect 55 785 98 802
rect 115 785 157 802
rect 174 785 216 802
rect 233 785 276 802
rect 293 785 335 802
rect 352 785 394 802
rect 411 785 439 802
rect 456 785 556 802
rect -63 762 -46 781
rect -46 745 -21 758
rect -63 741 -21 745
rect -4 741 46 758
rect 63 741 113 758
rect 130 741 180 758
rect 197 741 247 758
rect 264 741 315 758
rect 332 741 382 758
rect 399 741 425 758
rect 442 741 471 758
rect -63 721 -46 741
rect -63 702 -46 704
rect -159 685 -139 702
rect -122 685 -99 702
rect -82 685 -46 702
rect -29 685 -21 702
rect -4 685 38 702
rect 55 685 98 702
rect 115 685 157 702
rect 174 685 216 702
rect 233 685 276 702
rect 293 685 335 702
rect 352 685 394 702
rect 411 685 439 702
rect 456 685 505 702
rect -147 627 -130 685
rect -63 679 -46 685
rect -63 658 -46 662
rect -63 641 -21 658
rect -4 641 26 658
rect 43 641 64 658
rect 81 641 111 658
rect 128 641 158 658
rect 175 641 195 658
rect 212 641 243 658
rect 260 641 287 658
rect 304 641 327 658
rect 344 641 374 658
rect 391 641 433 658
rect 450 641 471 658
rect -63 636 -46 641
rect -147 592 -130 610
rect -147 549 -130 575
rect -147 507 -130 532
rect -147 464 -130 490
rect -147 422 -130 447
rect -147 379 -130 405
rect -147 337 -130 362
rect -147 294 -130 320
rect -147 252 -130 277
rect -147 209 -130 235
rect -147 160 -130 192
rect -147 135 -130 143
rect -103 627 -86 635
rect -103 592 -86 610
rect -103 549 -86 575
rect -103 507 -86 532
rect -103 464 -86 490
rect -103 422 -86 447
rect -103 379 -86 405
rect -103 337 -86 362
rect -103 294 -86 320
rect -103 252 -86 277
rect -103 209 -86 235
rect -103 160 -86 192
rect -103 110 -86 143
rect -63 594 -46 619
rect -29 585 -21 602
rect -4 585 38 602
rect 55 585 98 602
rect 115 585 157 602
rect 174 585 216 602
rect 233 585 276 602
rect 293 585 335 602
rect 352 585 385 602
rect 411 585 439 602
rect 456 585 471 602
rect -63 558 -46 577
rect -63 551 -21 558
rect -46 541 -21 551
rect -4 541 19 558
rect 36 541 75 558
rect 92 541 122 558
rect 139 541 171 558
rect 188 541 224 558
rect 241 541 268 558
rect 285 541 312 558
rect 329 541 364 558
rect 381 541 445 558
rect 462 541 471 558
rect -63 509 -46 534
rect -63 466 -46 492
rect -29 485 -21 502
rect -4 485 38 502
rect 55 485 98 502
rect 115 485 157 502
rect 174 485 216 502
rect 233 485 276 502
rect 293 485 335 502
rect 352 485 394 502
rect 411 485 439 502
rect 456 485 471 502
rect -46 449 -21 458
rect -63 441 -21 449
rect -4 441 32 458
rect 49 441 89 458
rect 106 441 134 458
rect 151 441 199 458
rect 216 441 237 458
rect 254 441 285 458
rect 302 441 329 458
rect 346 441 381 458
rect 398 441 442 458
rect 459 441 471 458
rect -63 424 -46 441
rect -63 381 -46 407
rect -29 385 -21 402
rect -4 385 38 402
rect 55 385 98 402
rect 115 385 157 402
rect 183 385 216 402
rect 233 385 276 402
rect 293 385 335 402
rect 352 385 394 402
rect 411 385 439 402
rect 456 385 471 402
rect -63 358 -46 364
rect -63 341 -21 358
rect -4 341 16 358
rect 33 341 75 358
rect 92 341 119 358
rect 136 341 171 358
rect 188 341 221 358
rect 238 341 267 358
rect 284 341 324 358
rect 341 341 363 358
rect 380 341 412 358
rect 429 341 446 358
rect 463 341 471 358
rect -63 339 -46 341
rect -63 296 -46 322
rect -29 285 -21 302
rect -4 285 38 302
rect 55 285 90 302
rect 115 285 157 302
rect 174 285 216 302
rect 233 285 276 302
rect 293 285 335 302
rect 352 285 394 302
rect 411 285 439 302
rect 456 285 471 302
rect -63 258 -46 279
rect -63 254 -21 258
rect -46 241 -21 254
rect -4 241 27 258
rect 44 241 86 258
rect 103 241 160 258
rect 177 241 234 258
rect 251 241 299 258
rect 316 241 363 258
rect 380 241 428 258
rect 445 241 471 258
rect -63 210 -46 237
rect -63 158 -46 193
rect -29 185 -21 202
rect 4 185 38 202
rect 55 185 98 202
rect 115 185 157 202
rect 174 185 216 202
rect 233 185 276 202
rect 293 185 335 202
rect 352 185 394 202
rect 411 185 439 202
rect 456 185 471 202
rect -46 141 -21 158
rect -4 141 36 158
rect 53 141 93 158
rect 110 141 150 158
rect 167 141 207 158
rect 224 141 264 158
rect 281 141 321 158
rect 338 141 378 158
rect 395 141 435 158
rect 452 141 460 158
rect 488 142 505 685
rect 477 125 505 142
rect 539 142 556 785
rect 577 571 594 819
rect 577 531 594 554
rect 577 491 594 514
rect 577 452 594 474
rect 577 412 594 435
rect 577 372 594 395
rect 577 332 594 355
rect 577 293 594 315
rect 577 253 594 276
rect 577 218 594 236
rect 577 184 594 201
rect 621 571 638 579
rect 621 531 638 554
rect 621 491 638 514
rect 621 452 638 474
rect 621 412 638 435
rect 621 372 638 395
rect 621 332 638 355
rect 621 293 638 315
rect 621 253 638 276
rect 621 218 638 236
rect 621 184 638 201
rect 615 167 621 184
rect 638 167 703 184
rect 577 159 594 167
rect 621 159 638 167
rect 539 125 594 142
rect -174 -171 -158 -154
rect -141 -171 -133 -154
rect -147 -209 -130 -201
rect -147 -244 -130 -226
rect -147 -279 -130 -261
rect -147 -314 -130 -296
rect -147 -348 -130 -331
rect -147 -383 -130 -365
rect -147 -418 -130 -400
rect -147 -453 -130 -435
rect -147 -488 -130 -470
rect -147 -523 -130 -505
rect -147 -558 -130 -540
rect -147 -592 -130 -575
rect -147 -627 -130 -609
rect -147 -676 -130 -644
rect -147 -751 -130 -693
rect -103 -209 -86 93
rect -23 63 -6 83
rect -23 25 -6 46
rect -23 0 -6 8
rect 21 100 38 108
rect 21 63 38 83
rect 21 23 38 46
rect 21 -25 38 6
rect 77 66 94 83
rect 77 25 94 49
rect 77 0 94 8
rect 121 100 138 108
rect 121 63 138 83
rect 121 23 138 46
rect 121 -25 138 6
rect 177 66 194 83
rect 177 25 194 49
rect 177 0 194 8
rect 221 100 238 108
rect 221 63 238 83
rect 221 23 238 46
rect 221 -25 238 6
rect 277 66 294 83
rect 277 25 294 49
rect 277 0 294 8
rect 321 100 338 108
rect 321 63 338 83
rect 321 23 338 46
rect 321 -25 338 6
rect 377 66 394 83
rect 377 25 394 49
rect 377 0 394 8
rect 421 100 438 108
rect 421 63 438 83
rect 421 23 438 46
rect 421 -25 438 6
rect 477 100 494 125
rect 477 66 494 83
rect 477 25 494 49
rect 477 0 494 8
rect 521 100 538 108
rect 521 66 538 83
rect 521 23 538 49
rect 521 -25 538 6
rect 577 100 594 125
rect 577 66 594 83
rect 577 25 594 49
rect 577 0 594 8
rect 621 100 638 108
rect 621 66 638 83
rect 621 23 638 49
rect 621 -24 638 6
rect 686 -24 703 167
rect -4 -42 4 -25
rect 21 -42 79 -25
rect 96 -42 104 -25
rect 121 -42 179 -25
rect 196 -42 204 -25
rect 221 -42 279 -25
rect 296 -42 304 -25
rect 321 -42 379 -25
rect 396 -42 404 -25
rect 421 -42 479 -25
rect 496 -42 504 -25
rect 521 -42 579 -25
rect 596 -42 604 -25
rect 621 -41 636 -24
rect 661 -41 669 -24
rect 686 -41 721 -24
rect -23 -74 -6 -66
rect -23 -111 -6 -91
rect -23 -149 -6 -128
rect -23 -207 -6 -166
rect 21 -72 38 -42
rect 21 -111 38 -89
rect 21 -149 38 -128
rect 21 -174 38 -166
rect 77 -74 94 -66
rect 77 -111 94 -91
rect 77 -149 94 -128
rect 121 -72 138 -42
rect 121 -112 138 -89
rect 121 -149 138 -129
rect 121 -174 138 -166
rect 177 -74 194 -66
rect 177 -111 194 -91
rect 177 -149 194 -128
rect 221 -72 238 -42
rect 221 -112 238 -89
rect 221 -149 238 -129
rect 221 -174 238 -166
rect 277 -74 294 -66
rect 277 -111 294 -91
rect 277 -149 294 -128
rect 321 -72 338 -42
rect 321 -111 338 -89
rect 321 -149 338 -128
rect 321 -174 338 -166
rect 377 -74 394 -66
rect 377 -111 394 -91
rect 377 -149 394 -128
rect 421 -72 438 -42
rect 421 -111 438 -89
rect 421 -149 438 -128
rect 421 -174 438 -166
rect 477 -74 494 -66
rect 477 -111 494 -91
rect 477 -149 494 -128
rect 477 -191 494 -166
rect 521 -74 538 -42
rect 521 -111 538 -91
rect 521 -149 538 -128
rect 521 -174 538 -166
rect 577 -74 594 -66
rect 577 -111 594 -91
rect 577 -149 594 -128
rect 577 -191 594 -166
rect 621 -74 638 -41
rect 621 -111 638 -91
rect 621 -149 638 -128
rect 621 -174 638 -166
rect -29 -224 -21 -207
rect -4 -224 56 -207
rect 73 -224 132 -207
rect 149 -224 209 -207
rect 226 -224 286 -207
rect 303 -224 362 -207
rect 379 -224 435 -207
rect 452 -224 460 -207
rect 477 -208 505 -191
rect -103 -244 -86 -226
rect -103 -279 -86 -261
rect -67 -249 -42 -243
rect -67 -263 -63 -249
rect -103 -314 -86 -296
rect -103 -348 -86 -331
rect -103 -383 -86 -365
rect -103 -418 -86 -400
rect -103 -453 -86 -435
rect -103 -488 -86 -470
rect -103 -523 -86 -505
rect -103 -558 -86 -540
rect -103 -592 -86 -575
rect -103 -627 -86 -609
rect -103 -676 -86 -644
rect -103 -701 -86 -693
rect -46 -251 -42 -249
rect -46 -266 -21 -251
rect -63 -268 -21 -266
rect -4 -268 24 -251
rect 41 -268 69 -251
rect 86 -268 113 -251
rect 130 -268 158 -251
rect 175 -268 203 -251
rect 220 -268 248 -251
rect 265 -268 293 -251
rect 310 -268 338 -251
rect 355 -268 383 -251
rect 400 -268 427 -251
rect 444 -268 471 -251
rect -63 -295 -46 -268
rect -63 -341 -46 -312
rect -29 -324 -21 -307
rect -4 -324 24 -307
rect 41 -324 69 -307
rect 94 -324 114 -307
rect 131 -324 159 -307
rect 176 -324 204 -307
rect 221 -324 248 -307
rect 265 -324 293 -307
rect 310 -324 338 -307
rect 355 -324 383 -307
rect 400 -324 428 -307
rect 445 -324 471 -307
rect -46 -358 -21 -351
rect -63 -368 -21 -358
rect -4 -368 24 -351
rect 41 -368 69 -351
rect 86 -368 113 -351
rect 130 -368 158 -351
rect 175 -368 203 -351
rect 220 -368 248 -351
rect 265 -368 293 -351
rect 310 -368 338 -351
rect 355 -368 383 -351
rect 400 -368 427 -351
rect 444 -368 471 -351
rect -63 -388 -46 -368
rect -63 -434 -46 -405
rect -29 -424 -21 -407
rect -4 -424 24 -407
rect 41 -424 69 -407
rect 86 -424 114 -407
rect 131 -424 170 -407
rect 196 -424 209 -407
rect 226 -424 248 -407
rect 265 -424 288 -407
rect 305 -424 327 -407
rect 344 -424 366 -407
rect 383 -424 405 -407
rect 422 -424 444 -407
rect 461 -424 471 -407
rect -63 -468 -21 -451
rect -4 -468 18 -451
rect 35 -468 58 -451
rect 75 -468 97 -451
rect 114 -468 136 -451
rect 153 -468 175 -451
rect 192 -468 214 -451
rect 231 -468 254 -451
rect 271 -468 293 -451
rect 310 -468 332 -451
rect 349 -468 371 -451
rect 388 -468 411 -451
rect 428 -468 445 -451
rect 462 -468 471 -451
rect -63 -480 -46 -468
rect -63 -527 -46 -497
rect -29 -524 -21 -507
rect -4 -524 18 -507
rect 35 -524 58 -507
rect 75 -524 97 -507
rect 114 -524 136 -507
rect 153 -524 175 -507
rect 192 -524 214 -507
rect 231 -524 254 -507
rect 271 -524 278 -507
rect 305 -524 327 -507
rect 344 -524 366 -507
rect 383 -524 406 -507
rect 423 -524 445 -507
rect 462 -524 471 -507
rect -63 -551 -46 -544
rect -63 -568 -21 -551
rect -4 -568 24 -551
rect 41 -568 69 -551
rect 86 -568 113 -551
rect 130 -568 158 -551
rect 175 -568 203 -551
rect 220 -568 248 -551
rect 265 -568 293 -551
rect 310 -568 338 -551
rect 355 -568 383 -551
rect 400 -568 427 -551
rect 444 -568 471 -551
rect -63 -573 -46 -568
rect -63 -619 -46 -590
rect -29 -624 -21 -607
rect -4 -624 24 -607
rect 41 -624 69 -607
rect 86 -624 114 -607
rect 131 -624 158 -607
rect 175 -624 203 -607
rect 220 -624 248 -607
rect 265 -624 293 -607
rect 310 -624 338 -607
rect 355 -624 378 -607
rect 400 -624 428 -607
rect 445 -624 471 -607
rect -63 -651 -46 -636
rect -63 -666 -21 -651
rect -46 -668 -21 -666
rect -4 -668 29 -651
rect 46 -668 80 -651
rect 97 -668 130 -651
rect 147 -668 181 -651
rect 198 -668 231 -651
rect 248 -668 282 -651
rect 299 -668 332 -651
rect 349 -668 383 -651
rect 400 -668 428 -651
rect 445 -668 471 -651
rect -63 -712 -46 -683
rect 488 -707 505 -208
rect -29 -724 -21 -707
rect -4 -724 24 -707
rect 41 -724 69 -707
rect 86 -724 114 -707
rect 131 -724 158 -707
rect 175 -724 203 -707
rect 220 -724 248 -707
rect 265 -724 293 -707
rect 310 -724 338 -707
rect 355 -724 383 -707
rect 400 -724 428 -707
rect 445 -724 505 -707
rect 522 -208 594 -191
rect -63 -751 -46 -729
rect -159 -768 -139 -751
rect -122 -768 -99 -751
rect -82 -758 -21 -751
rect -82 -768 -63 -758
rect -46 -768 -21 -758
rect -4 -768 24 -751
rect 41 -768 69 -751
rect 86 -768 113 -751
rect 130 -768 158 -751
rect 175 -768 203 -751
rect 220 -768 248 -751
rect 265 -768 293 -751
rect 310 -768 338 -751
rect 355 -768 373 -751
rect 390 -768 427 -751
rect 444 -768 471 -751
rect -63 -805 -46 -775
rect 522 -807 539 -208
rect -63 -851 -46 -822
rect -29 -824 -21 -807
rect -4 -824 24 -807
rect 41 -824 69 -807
rect 86 -824 113 -807
rect 130 -824 158 -807
rect 175 -824 203 -807
rect 220 -824 248 -807
rect 265 -824 293 -807
rect 310 -824 338 -807
rect 355 -824 383 -807
rect 400 -824 427 -807
rect 444 -824 539 -807
rect 577 -233 594 -225
rect 621 -233 638 -225
rect 686 -233 703 -41
rect 615 -250 621 -233
rect 638 -250 703 -233
rect 577 -271 594 -250
rect 577 -308 594 -288
rect 577 -851 594 -325
rect 621 -271 638 -250
rect 621 -308 638 -288
rect 621 -333 638 -325
rect -46 -868 -21 -851
rect -4 -868 24 -851
rect 41 -868 63 -851
rect 80 -868 102 -851
rect 119 -868 147 -851
rect 164 -868 192 -851
rect 209 -868 237 -851
rect 254 -868 282 -851
rect 299 -868 327 -851
rect 344 -868 371 -851
rect 388 -868 416 -851
rect 433 -868 450 -851
rect 467 -868 594 -851
rect -63 -885 -46 -868
rect -21 -885 -4 -868
rect 24 -885 41 -868
rect 63 -885 80 -868
rect 102 -885 119 -868
rect 147 -885 164 -868
rect 192 -885 209 -868
rect 237 -885 254 -868
rect 282 -885 299 -868
rect 327 -885 344 -868
rect 371 -885 388 -868
rect 416 -885 433 -868
rect 450 -885 467 -868
rect -63 -889 676 -885
rect -63 -890 653 -889
rect -63 -907 -55 -890
rect -38 -907 -6 -890
rect 11 -907 55 -890
rect 72 -907 117 -890
rect 134 -907 178 -890
rect 195 -907 240 -890
rect 257 -907 301 -890
rect 318 -907 363 -890
rect 380 -907 424 -890
rect 441 -907 486 -890
rect 503 -907 547 -890
rect 564 -907 609 -890
rect 626 -906 653 -890
rect 670 -906 676 -889
rect 626 -907 676 -906
rect -63 -910 676 -907
<< viali >>
rect -55 823 -38 840
rect -18 823 -1 840
rect 26 823 43 840
rect 71 823 88 840
rect 115 823 132 840
rect 159 823 176 840
rect 204 823 221 840
rect 248 823 265 840
rect 292 823 309 840
rect 336 823 353 840
rect 381 823 398 840
rect 425 823 442 840
rect 469 823 486 840
rect 514 823 531 840
rect 558 823 575 840
rect 602 823 619 840
rect 647 823 664 840
rect -63 781 -46 798
rect -63 745 -46 762
rect -63 704 -46 721
rect -139 685 -122 702
rect -99 685 -82 702
rect -63 662 -46 679
rect -63 619 -46 636
rect -63 577 -46 594
rect 385 585 394 602
rect 394 585 402 602
rect -63 534 -46 551
rect -63 492 -46 509
rect 276 485 293 502
rect -63 449 -46 466
rect -63 407 -46 424
rect 166 385 174 402
rect 174 385 183 402
rect -63 364 -46 381
rect -63 322 -46 339
rect -63 279 -46 296
rect 90 285 98 302
rect 98 285 107 302
rect -63 237 -46 254
rect -63 193 -46 210
rect -13 185 -4 202
rect -4 185 4 202
rect -63 141 -46 158
rect -23 100 -6 108
rect -23 91 -6 100
rect 77 100 94 108
rect 77 91 94 100
rect 177 100 194 108
rect 177 91 194 100
rect 277 100 294 108
rect 277 91 294 100
rect 377 100 394 108
rect 377 91 394 100
rect -29 -42 -21 -25
rect -21 -42 -12 -25
rect 636 -41 644 -24
rect 644 -41 653 -24
rect 77 -166 94 -157
rect 77 -174 94 -166
rect 177 -166 194 -157
rect 177 -174 194 -166
rect 277 -166 294 -157
rect 277 -174 294 -166
rect 377 -166 394 -157
rect 377 -174 394 -166
rect -63 -266 -46 -249
rect -63 -312 -46 -295
rect 77 -324 86 -307
rect 86 -324 94 -307
rect -63 -358 -46 -341
rect -63 -405 -46 -388
rect 179 -424 187 -407
rect 187 -424 196 -407
rect -63 -451 -46 -434
rect -63 -497 -46 -480
rect 278 -524 288 -507
rect 288 -524 295 -507
rect -63 -544 -46 -527
rect -63 -590 -46 -573
rect -63 -636 -46 -619
rect 378 -624 383 -607
rect 383 -624 395 -607
rect -63 -683 -46 -666
rect -63 -729 -46 -712
rect -139 -768 -122 -751
rect -99 -768 -82 -751
rect -63 -775 -46 -758
rect -63 -822 -46 -805
rect -63 -868 -46 -851
rect -55 -907 -38 -890
rect -6 -907 11 -890
rect 55 -907 72 -890
rect 117 -907 134 -890
rect 178 -907 195 -890
rect 240 -907 257 -890
rect 301 -907 318 -890
rect 363 -907 380 -890
rect 424 -907 441 -890
rect 486 -907 503 -890
rect 547 -907 564 -890
rect 609 -907 626 -890
rect 653 -906 670 -889
<< metal1 >>
rect -67 840 670 844
rect -67 823 -55 840
rect -38 823 -18 840
rect -1 823 26 840
rect 43 823 71 840
rect 88 823 115 840
rect 132 823 159 840
rect 176 823 204 840
rect 221 823 248 840
rect 265 823 292 840
rect 309 823 336 840
rect 353 823 381 840
rect 398 823 425 840
rect 442 823 469 840
rect 486 823 514 840
rect 531 823 558 840
rect 575 823 602 840
rect 619 823 647 840
rect 664 823 670 840
rect -67 819 670 823
rect -67 798 -42 819
rect -67 781 -63 798
rect -46 781 -42 798
rect -67 762 -42 781
rect -67 745 -63 762
rect -46 745 -42 762
rect -67 721 -42 745
rect -67 706 -63 721
rect -147 704 -63 706
rect -46 704 -42 721
rect -147 702 -42 704
rect -147 685 -139 702
rect -122 685 -99 702
rect -82 685 -42 702
rect -147 681 -42 685
rect -67 679 -42 681
rect -67 662 -63 679
rect -46 662 -42 679
rect -67 636 -42 662
rect -67 619 -63 636
rect -46 619 -42 636
rect -67 594 -42 619
rect -67 577 -63 594
rect -46 577 -42 594
rect -67 551 -42 577
rect -67 534 -63 551
rect -46 534 -42 551
rect -67 509 -42 534
rect -67 492 -63 509
rect -46 492 -42 509
rect 371 602 411 608
rect 371 585 385 602
rect 402 585 411 602
rect 371 579 411 585
rect -67 466 -42 492
rect -67 449 -63 466
rect -46 449 -42 466
rect -67 424 -42 449
rect -67 407 -63 424
rect -46 407 -42 424
rect 271 502 300 508
rect 271 485 276 502
rect 293 485 300 502
rect -67 381 -42 407
rect -67 364 -63 381
rect -46 364 -42 381
rect 157 402 200 408
rect 157 385 166 402
rect 183 385 200 402
rect 157 379 200 385
rect -67 339 -42 364
rect -67 322 -63 339
rect -46 322 -42 339
rect -67 296 -42 322
rect -67 279 -63 296
rect -46 279 -42 296
rect -67 254 -42 279
rect -67 237 -63 254
rect -46 237 -42 254
rect -67 210 -42 237
rect -67 193 -63 210
rect -46 193 -42 210
rect 71 302 115 308
rect 71 285 90 302
rect 107 285 115 302
rect 71 279 115 285
rect -67 158 -42 193
rect -67 141 -63 158
rect -46 141 -42 158
rect -67 135 -42 141
rect -28 202 11 208
rect -28 185 -13 202
rect 4 185 11 202
rect -28 179 11 185
rect -28 108 -1 179
rect -28 91 -23 108
rect -6 91 -1 108
rect -28 83 -1 91
rect 71 108 100 279
rect 71 91 77 108
rect 94 91 100 108
rect 71 83 100 91
rect 171 108 200 379
rect 171 91 177 108
rect 194 91 200 108
rect 171 83 200 91
rect 271 108 300 485
rect 271 91 277 108
rect 294 91 300 108
rect 271 83 300 91
rect 371 108 400 579
rect 371 91 377 108
rect 394 91 400 108
rect 371 83 400 91
rect -47 -24 662 -18
rect -47 -25 636 -24
rect -47 -42 -29 -25
rect -12 -41 636 -25
rect 653 -41 662 -24
rect -12 -42 662 -41
rect -47 -49 662 -42
rect 71 -157 100 -149
rect 71 -174 77 -157
rect 94 -174 100 -157
rect -67 -249 -42 -243
rect -67 -266 -63 -249
rect -46 -266 -42 -249
rect -67 -295 -42 -266
rect -67 -312 -63 -295
rect -46 -312 -42 -295
rect -67 -341 -42 -312
rect 71 -307 100 -174
rect 71 -324 77 -307
rect 94 -324 100 -307
rect 71 -330 100 -324
rect 171 -157 200 -149
rect 171 -174 177 -157
rect 194 -174 200 -157
rect -67 -358 -63 -341
rect -46 -358 -42 -341
rect -67 -388 -42 -358
rect -67 -405 -63 -388
rect -46 -405 -42 -388
rect -67 -434 -42 -405
rect 171 -407 200 -174
rect 171 -424 179 -407
rect 196 -424 200 -407
rect 171 -430 200 -424
rect 271 -157 300 -149
rect 271 -174 277 -157
rect 294 -174 300 -157
rect -67 -451 -63 -434
rect -46 -451 -42 -434
rect -67 -480 -42 -451
rect -67 -497 -63 -480
rect -46 -497 -42 -480
rect -67 -527 -42 -497
rect -67 -544 -63 -527
rect -46 -544 -42 -527
rect 271 -507 300 -174
rect 271 -524 278 -507
rect 295 -524 300 -507
rect 271 -530 300 -524
rect 371 -157 400 -149
rect 371 -174 377 -157
rect 394 -174 400 -157
rect -67 -573 -42 -544
rect -67 -590 -63 -573
rect -46 -590 -42 -573
rect -67 -619 -42 -590
rect -67 -636 -63 -619
rect -46 -636 -42 -619
rect 371 -607 400 -174
rect 371 -624 378 -607
rect 395 -624 400 -607
rect 371 -630 400 -624
rect -67 -666 -42 -636
rect -67 -683 -63 -666
rect -46 -683 -42 -666
rect -67 -712 -42 -683
rect -67 -729 -63 -712
rect -46 -729 -42 -712
rect -67 -747 -42 -729
rect -147 -751 -42 -747
rect -147 -768 -139 -751
rect -122 -768 -99 -751
rect -82 -758 -42 -751
rect -82 -768 -63 -758
rect -147 -772 -63 -768
rect -67 -775 -63 -772
rect -46 -775 -42 -758
rect -67 -805 -42 -775
rect -67 -822 -63 -805
rect -46 -822 -42 -805
rect -67 -851 -42 -822
rect -67 -868 -63 -851
rect -46 -868 -42 -851
rect -67 -885 -42 -868
rect -67 -889 676 -885
rect -67 -890 653 -889
rect -67 -907 -55 -890
rect -38 -907 -6 -890
rect 11 -907 55 -890
rect 72 -907 117 -890
rect 134 -907 178 -890
rect 195 -907 240 -890
rect 257 -907 301 -890
rect 318 -907 363 -890
rect 380 -907 424 -890
rect 441 -907 486 -890
rect 503 -907 547 -890
rect 564 -907 609 -890
rect 626 -906 653 -890
rect 670 -906 676 -889
rect 626 -907 676 -906
rect -67 -910 676 -907
<< labels >>
rlabel locali -174 -171 -174 -154 3 in
port 1 e
rlabel locali -159 685 -159 702 1 vdd
port 3 n
rlabel locali -159 -768 -159 -751 1 gnd
port 4 n
rlabel locali 721 -41 721 -24 7 out
port 5 w
<< end >>
