*PLL
.include sky130nm.lib

xx1 Clk_Ref Clk_Out_by_8 up down pd
xx2 up down VCtrl cp

*Loop Filter
r1 VCtrl rc1 490
c1 rc1 0 355f
r2 rc1 rc2 490
c2 rc2 0 350f
r3 rc2 rc3 490
c3 rc3 0 345f

xx3 rc3 Clk_Out vco

xx4 Clk_Out Clk_Out_by_2 fd
xx5 Clk_Out_by_2 Clk_Out_by_4 fd
xx6 Clk_Out_by_4 Clk_Out_by_8 fd

v1 Clk_Ref 0 PULSE 0 1.8 0 6ps 6ps 40ns 80ns

.ic v(VCtrl) = 0
.ic v(Clk_Out_by_2) = 0
.ic v(Clk_Out_by_4) = 1.8
.ic v(Clk_Out_by_8) = 0
.control
tran 0.1ns 180us
plot v(Clk_Ref) v(Clk_Out_by_8) v(Clk_Out_by_4)+2 v(Clk_Out_by_2)+4 v(Clk_Out)+6 v(up)+8 v(down)+10 v(VCtrl)+12
.endc

*PFD
.subckt pd Clk1 Clk2 up down 
xm1 1 clk1 3 1 sky130_fd_pr__pfet_01v8 l=150n w=640n 
xm2 3 clk1 4 0 sky130_fd_pr__nfet_01v8 l=150n w=1800n
xm3 4 clk2 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 clk2 6 1 sky130_fd_pr__pfet_01v8 l=150n w=640n 
xm5 6 clk2 7 0 sky130_fd_pr__nfet_01v8 l=150n w=1800n
xm6 7 clk1 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm7 8 clk1 3 0 sky130_fd_pr__nfet_01v8 l=150n w=2400n 
xm8 clk1 clk1 8 1 sky130_fd_pr__pfet_01v8 l=150n w=640n

xm11 upb 8 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm12 upb 8 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm15 up upb 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm16 up upb 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
  
xm9 9 clk2 6 0 sky130_fd_pr__nfet_01v8 l=150n w=2400n
xm10 clk2 clk2 9 1 sky130_fd_pr__pfet_01v8 l=150n w=640n

xm13 downb 9 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm14 downb 9 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm17 down downb 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm18 down downb 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n


*output cap
*c1 up 0 6f
*c2 down 0 6f

v1 1 0 1.8
.ends pd


*CP
.subckt cp up down out
xm43 3 2 1 1 sky130_fd_pr__pfet_01v8 l=150n w=18u 
xm44 out downb 3 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm31 out up 7 0 sky130_fd_pr__nfet_01v8 l=150n w=420n
xm32 7 8 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4.8u

xm33 2 2 1 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm34 8 8 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm35 9 down 3 1 sky130_fd_pr__pfet_01v8 l=150n w=5400n 
xm36 9 9 0 0 sky130_fd_pr__nfet_01v8 l=150n w=420n

xm37 10 10 1 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm38 10 upb 7 0 sky130_fd_pr__nfet_01v8 l=150n w=5400n

xm39 1 down downb 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm40 0 down downb 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 

xm41 1 up upb 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm42 0 up upb 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 

*r1 out rc 200
*c1 rc 0 8f

v1 1 0 1.8
.ends cp


*VCO
.subckt vco in out
XM1 A A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM2 A in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM3 C A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM4 H in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM5 D A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM6 I in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM7 E A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM8 J in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM9 F A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM10 K in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM11 G A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM12 L in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM13 R A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM14 T in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM15 S A 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM16 U in 0 0 sky130_fd_pr__nfet_01v8 l=150n w=4200n

XM17 M Z C C sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM18 M Z H H sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM19 N M D D sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM20 N M I I sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM21 O N E E sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM22 O N J J sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM23 P O F F sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM24 P O K K sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM25 Q P G G sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM26 Q P L L sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM27 V Q R R sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM28 V Q T T sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM29 Z V S S sky130_fd_pr__pfet_01v8 l=150n w=1080n
XM30 Z V U U sky130_fd_pr__nfet_01v8 l=150n w=1080n

XM31 out Z 1 1 sky130_fd_pr__pfet_01v8 l=150n w=4200n
XM32 out Z 0 0 sky130_fd_pr__nfet_01v8 l=150n w=1080n

*c1 11 0 24f
v1 1 0 1.8
.ends vco


*FD
.subckt fd Clk 10

xm1 1 2 3 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm2 0 2 3 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 

xm3 3 Clkb 4 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm4 3 Clk 4 0 sky130_fd_pr__nfet_01v8 l=150n w=840n 

xm7 1 4 5 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm8 0 4 5 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 

xm9 5 Clk 6 1 sky130_fd_pr__pfet_01v8 l=150n w=420n 
xm10 5 Clkb 6 0 sky130_fd_pr__nfet_01v8 l=150n w=640n 

xm11 1 6 2 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm12 0 6 2 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 

xm13 1 Clk Clkb 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm14 0 Clk Clkb 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 

xm15 7 6 1 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
xm16 7 6 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm19 1 7 10 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm20 10 7 0 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 


*c1 7 0 18f
v1 1 0 1.8
.ends fd